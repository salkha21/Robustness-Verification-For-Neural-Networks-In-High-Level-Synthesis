module test_linear_tb;

    // Parameters
    parameter CLK_PERIOD = 10; // Clock period in nanoseconds

    // Inputs
    reg clk;
    reg rst;


    reg [11:0] p__arg0_0_0;
	reg [11:0] p__arg0_0_1;
	reg [11:0] p__arg0_0_10;
	reg [11:0] p__arg0_0_2;
	reg [11:0] p__arg0_0_3;
	reg [11:0] p__arg0_0_4;
	reg [11:0] p__arg0_0_5;
	reg [11:0] p__arg0_0_6;
	reg [11:0] p__arg0_0_7;
	reg [11:0] p__arg0_0_8;
	reg [11:0] p__arg0_0_9;
	reg [11:0] p___constant_11x11xf32_0_0;
	reg [11:0] p___constant_11x11xf32_0_1;
	reg [11:0] p___constant_11x11xf32_0_10;
	reg [11:0] p___constant_11x11xf32_0_2;
	reg [11:0] p___constant_11x11xf32_0_3;
	reg [11:0] p___constant_11x11xf32_0_4;
	reg [11:0] p___constant_11x11xf32_0_5;
	reg [11:0] p___constant_11x11xf32_0_6;
	reg [11:0] p___constant_11x11xf32_0_7;
	reg [11:0] p___constant_11x11xf32_0_8;
	reg [11:0] p___constant_11x11xf32_0_9;
	reg [11:0] p___constant_11x11xf32_10_0;
	reg [11:0] p___constant_11x11xf32_10_1;
	reg [11:0] p___constant_11x11xf32_10_10;
	reg [11:0] p___constant_11x11xf32_10_2;
	reg [11:0] p___constant_11x11xf32_10_3;
	reg [11:0] p___constant_11x11xf32_10_4;
	reg [11:0] p___constant_11x11xf32_10_5;
	reg [11:0] p___constant_11x11xf32_10_6;
	reg [11:0] p___constant_11x11xf32_10_7;
	reg [11:0] p___constant_11x11xf32_10_8;
	reg [11:0] p___constant_11x11xf32_10_9;
	reg [11:0] p___constant_11x11xf32_1_0;
	reg [11:0] p___constant_11x11xf32_1_1;
	reg [11:0] p___constant_11x11xf32_1_10;
	reg [11:0] p___constant_11x11xf32_1_2;
	reg [11:0] p___constant_11x11xf32_1_3;
	reg [11:0] p___constant_11x11xf32_1_4;
	reg [11:0] p___constant_11x11xf32_1_5;
	reg [11:0] p___constant_11x11xf32_1_6;
	reg [11:0] p___constant_11x11xf32_1_7;
	reg [11:0] p___constant_11x11xf32_1_8;
	reg [11:0] p___constant_11x11xf32_1_9;
	reg [11:0] p___constant_11x11xf32_2_0;
	reg [11:0] p___constant_11x11xf32_2_1;
	reg [11:0] p___constant_11x11xf32_2_10;
	reg [11:0] p___constant_11x11xf32_2_2;
	reg [11:0] p___constant_11x11xf32_2_3;
	reg [11:0] p___constant_11x11xf32_2_4;
	reg [11:0] p___constant_11x11xf32_2_5;
	reg [11:0] p___constant_11x11xf32_2_6;
	reg [11:0] p___constant_11x11xf32_2_7;
	reg [11:0] p___constant_11x11xf32_2_8;
	reg [11:0] p___constant_11x11xf32_2_9;
	reg [11:0] p___constant_11x11xf32_3_0;
	reg [11:0] p___constant_11x11xf32_3_1;
	reg [11:0] p___constant_11x11xf32_3_10;
	reg [11:0] p___constant_11x11xf32_3_2;
	reg [11:0] p___constant_11x11xf32_3_3;
	reg [11:0] p___constant_11x11xf32_3_4;
	reg [11:0] p___constant_11x11xf32_3_5;
	reg [11:0] p___constant_11x11xf32_3_6;
	reg [11:0] p___constant_11x11xf32_3_7;
	reg [11:0] p___constant_11x11xf32_3_8;
	reg [11:0] p___constant_11x11xf32_3_9;
	reg [11:0] p___constant_11x11xf32_4_0;
	reg [11:0] p___constant_11x11xf32_4_1;
	reg [11:0] p___constant_11x11xf32_4_10;
	reg [11:0] p___constant_11x11xf32_4_2;
	reg [11:0] p___constant_11x11xf32_4_3;
	reg [11:0] p___constant_11x11xf32_4_4;
	reg [11:0] p___constant_11x11xf32_4_5;
	reg [11:0] p___constant_11x11xf32_4_6;
	reg [11:0] p___constant_11x11xf32_4_7;
	reg [11:0] p___constant_11x11xf32_4_8;
	reg [11:0] p___constant_11x11xf32_4_9;
	reg [11:0] p___constant_11x11xf32_5_0;
	reg [11:0] p___constant_11x11xf32_5_1;
	reg [11:0] p___constant_11x11xf32_5_10;
	reg [11:0] p___constant_11x11xf32_5_2;
	reg [11:0] p___constant_11x11xf32_5_3;
	reg [11:0] p___constant_11x11xf32_5_4;
	reg [11:0] p___constant_11x11xf32_5_5;
	reg [11:0] p___constant_11x11xf32_5_6;
	reg [11:0] p___constant_11x11xf32_5_7;
	reg [11:0] p___constant_11x11xf32_5_8;
	reg [11:0] p___constant_11x11xf32_5_9;
	reg [11:0] p___constant_11x11xf32_6_0;
	reg [11:0] p___constant_11x11xf32_6_1;
	reg [11:0] p___constant_11x11xf32_6_10;
	reg [11:0] p___constant_11x11xf32_6_2;
	reg [11:0] p___constant_11x11xf32_6_3;
	reg [11:0] p___constant_11x11xf32_6_4;
	reg [11:0] p___constant_11x11xf32_6_5;
	reg [11:0] p___constant_11x11xf32_6_6;
	reg [11:0] p___constant_11x11xf32_6_7;
	reg [11:0] p___constant_11x11xf32_6_8;
	reg [11:0] p___constant_11x11xf32_6_9;
	reg [11:0] p___constant_11x11xf32_7_0;
	reg [11:0] p___constant_11x11xf32_7_1;
	reg [11:0] p___constant_11x11xf32_7_10;
	reg [11:0] p___constant_11x11xf32_7_2;
	reg [11:0] p___constant_11x11xf32_7_3;
	reg [11:0] p___constant_11x11xf32_7_4;
	reg [11:0] p___constant_11x11xf32_7_5;
	reg [11:0] p___constant_11x11xf32_7_6;
	reg [11:0] p___constant_11x11xf32_7_7;
	reg [11:0] p___constant_11x11xf32_7_8;
	reg [11:0] p___constant_11x11xf32_7_9;
	reg [11:0] p___constant_11x11xf32_8_0;
	reg [11:0] p___constant_11x11xf32_8_1;
	reg [11:0] p___constant_11x11xf32_8_10;
	reg [11:0] p___constant_11x11xf32_8_2;
	reg [11:0] p___constant_11x11xf32_8_3;
	reg [11:0] p___constant_11x11xf32_8_4;
	reg [11:0] p___constant_11x11xf32_8_5;
	reg [11:0] p___constant_11x11xf32_8_6;
	reg [11:0] p___constant_11x11xf32_8_7;
	reg [11:0] p___constant_11x11xf32_8_8;
	reg [11:0] p___constant_11x11xf32_8_9;
	reg [11:0] p___constant_11x11xf32_9_0;
	reg [11:0] p___constant_11x11xf32_9_1;
	reg [11:0] p___constant_11x11xf32_9_10;
	reg [11:0] p___constant_11x11xf32_9_2;
	reg [11:0] p___constant_11x11xf32_9_3;
	reg [11:0] p___constant_11x11xf32_9_4;
	reg [11:0] p___constant_11x11xf32_9_5;
	reg [11:0] p___constant_11x11xf32_9_6;
	reg [11:0] p___constant_11x11xf32_9_7;
	reg [11:0] p___constant_11x11xf32_9_8;
	reg [11:0] p___constant_11x11xf32_9_9;
	reg [11:0] p___constant_11xf32_0;
	reg [11:0] p___constant_11xf32_1;
	reg [11:0] p___constant_11xf32_10;
	reg [11:0] p___constant_11xf32_2;
	reg [11:0] p___constant_11xf32_3;
	reg [11:0] p___constant_11xf32_4;
	reg [11:0] p___constant_11xf32_5;
	reg [11:0] p___constant_11xf32_6;
	reg [11:0] p___constant_11xf32_7;
	reg [11:0] p___constant_11xf32_8;
	reg [11:0] p___constant_11xf32_9;
	wire [11:0] output_p_val_313;

    linear uut(
        .clk(clk),
        .rst(rst),
        .p__arg0_0_0(p__arg0_0_0),
        .p__arg0_0_1(p__arg0_0_1),
        .p__arg0_0_10(p__arg0_0_10),
        .p__arg0_0_2(p__arg0_0_2),
        .p__arg0_0_3(p__arg0_0_3),
        .p__arg0_0_4(p__arg0_0_4),
        .p__arg0_0_5(p__arg0_0_5),
        .p__arg0_0_6(p__arg0_0_6),
        .p__arg0_0_7(p__arg0_0_7),
        .p__arg0_0_8(p__arg0_0_8),
        .p__arg0_0_9(p__arg0_0_9),
        .p___constant_11x11xf32_0_0(p___constant_11x11xf32_0_0),
        .p___constant_11x11xf32_0_1(p___constant_11x11xf32_0_1),
        .p___constant_11x11xf32_0_10(p___constant_11x11xf32_0_10),
        .p___constant_11x11xf32_0_2(p___constant_11x11xf32_0_2),
        .p___constant_11x11xf32_0_3(p___constant_11x11xf32_0_3),
        .p___constant_11x11xf32_0_4(p___constant_11x11xf32_0_4),
        .p___constant_11x11xf32_0_5(p___constant_11x11xf32_0_5),
        .p___constant_11x11xf32_0_6(p___constant_11x11xf32_0_6),
        .p___constant_11x11xf32_0_7(p___constant_11x11xf32_0_7),
        .p___constant_11x11xf32_0_8(p___constant_11x11xf32_0_8),
        .p___constant_11x11xf32_0_9(p___constant_11x11xf32_0_9),
        .p___constant_11x11xf32_10_0(p___constant_11x11xf32_10_0),
        .p___constant_11x11xf32_10_1(p___constant_11x11xf32_10_1),
        .p___constant_11x11xf32_10_10(p___constant_11x11xf32_10_10),
        .p___constant_11x11xf32_10_2(p___constant_11x11xf32_10_2),
        .p___constant_11x11xf32_10_3(p___constant_11x11xf32_10_3),
        .p___constant_11x11xf32_10_4(p___constant_11x11xf32_10_4),
        .p___constant_11x11xf32_10_5(p___constant_11x11xf32_10_5),
        .p___constant_11x11xf32_10_6(p___constant_11x11xf32_10_6),
        .p___constant_11x11xf32_10_7(p___constant_11x11xf32_10_7),
        .p___constant_11x11xf32_10_8(p___constant_11x11xf32_10_8),
        .p___constant_11x11xf32_10_9(p___constant_11x11xf32_10_9),
        .p___constant_11x11xf32_1_0(p___constant_11x11xf32_1_0),
        .p___constant_11x11xf32_1_1(p___constant_11x11xf32_1_1),
        .p___constant_11x11xf32_1_10(p___constant_11x11xf32_1_10),
        .p___constant_11x11xf32_1_2(p___constant_11x11xf32_1_2),
        .p___constant_11x11xf32_1_3(p___constant_11x11xf32_1_3),
        .p___constant_11x11xf32_1_4(p___constant_11x11xf32_1_4),
        .p___constant_11x11xf32_1_5(p___constant_11x11xf32_1_5),
        .p___constant_11x11xf32_1_6(p___constant_11x11xf32_1_6),
        .p___constant_11x11xf32_1_7(p___constant_11x11xf32_1_7),
        .p___constant_11x11xf32_1_8(p___constant_11x11xf32_1_8),
        .p___constant_11x11xf32_1_9(p___constant_11x11xf32_1_9),
        .p___constant_11x11xf32_2_0(p___constant_11x11xf32_2_0),
        .p___constant_11x11xf32_2_1(p___constant_11x11xf32_2_1),
        .p___constant_11x11xf32_2_10(p___constant_11x11xf32_2_10),
        .p___constant_11x11xf32_2_2(p___constant_11x11xf32_2_2),
        .p___constant_11x11xf32_2_3(p___constant_11x11xf32_2_3),
        .p___constant_11x11xf32_2_4(p___constant_11x11xf32_2_4),
        .p___constant_11x11xf32_2_5(p___constant_11x11xf32_2_5),
        .p___constant_11x11xf32_2_6(p___constant_11x11xf32_2_6),
        .p___constant_11x11xf32_2_7(p___constant_11x11xf32_2_7),
        .p___constant_11x11xf32_2_8(p___constant_11x11xf32_2_8),
        .p___constant_11x11xf32_2_9(p___constant_11x11xf32_2_9),
        .p___constant_11x11xf32_3_0(p___constant_11x11xf32_3_0),
        .p___constant_11x11xf32_3_1(p___constant_11x11xf32_3_1),
        .p___constant_11x11xf32_3_10(p___constant_11x11xf32_3_10),
        .p___constant_11x11xf32_3_2(p___constant_11x11xf32_3_2),
        .p___constant_11x11xf32_3_3(p___constant_11x11xf32_3_3),
        .p___constant_11x11xf32_3_4(p___constant_11x11xf32_3_4),
        .p___constant_11x11xf32_3_5(p___constant_11x11xf32_3_5),
        .p___constant_11x11xf32_3_6(p___constant_11x11xf32_3_6),
        .p___constant_11x11xf32_3_7(p___constant_11x11xf32_3_7),
        .p___constant_11x11xf32_3_8(p___constant_11x11xf32_3_8),
        .p___constant_11x11xf32_3_9(p___constant_11x11xf32_3_9),
        .p___constant_11x11xf32_4_0(p___constant_11x11xf32_4_0),
        .p___constant_11x11xf32_4_1(p___constant_11x11xf32_4_1),
        .p___constant_11x11xf32_4_10(p___constant_11x11xf32_4_10),
        .p___constant_11x11xf32_4_2(p___constant_11x11xf32_4_2),
        .p___constant_11x11xf32_4_3(p___constant_11x11xf32_4_3),
        .p___constant_11x11xf32_4_4(p___constant_11x11xf32_4_4),
        .p___constant_11x11xf32_4_5(p___constant_11x11xf32_4_5),
        .p___constant_11x11xf32_4_6(p___constant_11x11xf32_4_6),
        .p___constant_11x11xf32_4_7(p___constant_11x11xf32_4_7),
        .p___constant_11x11xf32_4_8(p___constant_11x11xf32_4_8),
        .p___constant_11x11xf32_4_9(p___constant_11x11xf32_4_9),
        .p___constant_11x11xf32_5_0(p___constant_11x11xf32_5_0),
        .p___constant_11x11xf32_5_1(p___constant_11x11xf32_5_1),
        .p___constant_11x11xf32_5_10(p___constant_11x11xf32_5_10),
        .p___constant_11x11xf32_5_2(p___constant_11x11xf32_5_2),
        .p___constant_11x11xf32_5_3(p___constant_11x11xf32_5_3),
        .p___constant_11x11xf32_5_4(p___constant_11x11xf32_5_4),
        .p___constant_11x11xf32_5_5(p___constant_11x11xf32_5_5),
        .p___constant_11x11xf32_5_6(p___constant_11x11xf32_5_6),
        .p___constant_11x11xf32_5_7(p___constant_11x11xf32_5_7),
        .p___constant_11x11xf32_5_8(p___constant_11x11xf32_5_8),
        .p___constant_11x11xf32_5_9(p___constant_11x11xf32_5_9),
        .p___constant_11x11xf32_6_0(p___constant_11x11xf32_6_0),
        .p___constant_11x11xf32_6_1(p___constant_11x11xf32_6_1),
        .p___constant_11x11xf32_6_10(p___constant_11x11xf32_6_10),
        .p___constant_11x11xf32_6_2(p___constant_11x11xf32_6_2),
        .p___constant_11x11xf32_6_3(p___constant_11x11xf32_6_3),
        .p___constant_11x11xf32_6_4(p___constant_11x11xf32_6_4),
        .p___constant_11x11xf32_6_5(p___constant_11x11xf32_6_5),
        .p___constant_11x11xf32_6_6(p___constant_11x11xf32_6_6),
        .p___constant_11x11xf32_6_7(p___constant_11x11xf32_6_7),
        .p___constant_11x11xf32_6_8(p___constant_11x11xf32_6_8),
        .p___constant_11x11xf32_6_9(p___constant_11x11xf32_6_9),
        .p___constant_11x11xf32_7_0(p___constant_11x11xf32_7_0),
        .p___constant_11x11xf32_7_1(p___constant_11x11xf32_7_1),
        .p___constant_11x11xf32_7_10(p___constant_11x11xf32_7_10),
        .p___constant_11x11xf32_7_2(p___constant_11x11xf32_7_2),
        .p___constant_11x11xf32_7_3(p___constant_11x11xf32_7_3),
        .p___constant_11x11xf32_7_4(p___constant_11x11xf32_7_4),
        .p___constant_11x11xf32_7_5(p___constant_11x11xf32_7_5),
        .p___constant_11x11xf32_7_6(p___constant_11x11xf32_7_6),
        .p___constant_11x11xf32_7_7(p___constant_11x11xf32_7_7),
        .p___constant_11x11xf32_7_8(p___constant_11x11xf32_7_8),
        .p___constant_11x11xf32_7_9(p___constant_11x11xf32_7_9),
        .p___constant_11x11xf32_8_0(p___constant_11x11xf32_8_0),
        .p___constant_11x11xf32_8_1(p___constant_11x11xf32_8_1),
        .p___constant_11x11xf32_8_10(p___constant_11x11xf32_8_10),
        .p___constant_11x11xf32_8_2(p___constant_11x11xf32_8_2),
        .p___constant_11x11xf32_8_3(p___constant_11x11xf32_8_3),
        .p___constant_11x11xf32_8_4(p___constant_11x11xf32_8_4),
        .p___constant_11x11xf32_8_5(p___constant_11x11xf32_8_5),
        .p___constant_11x11xf32_8_6(p___constant_11x11xf32_8_6),
        .p___constant_11x11xf32_8_7(p___constant_11x11xf32_8_7),
        .p___constant_11x11xf32_8_8(p___constant_11x11xf32_8_8),
        .p___constant_11x11xf32_8_9(p___constant_11x11xf32_8_9),
        .p___constant_11x11xf32_9_0(p___constant_11x11xf32_9_0),
        .p___constant_11x11xf32_9_1(p___constant_11x11xf32_9_1),
        .p___constant_11x11xf32_9_10(p___constant_11x11xf32_9_10),
        .p___constant_11x11xf32_9_2(p___constant_11x11xf32_9_2),
        .p___constant_11x11xf32_9_3(p___constant_11x11xf32_9_3),
        .p___constant_11x11xf32_9_4(p___constant_11x11xf32_9_4),
        .p___constant_11x11xf32_9_5(p___constant_11x11xf32_9_5),
        .p___constant_11x11xf32_9_6(p___constant_11x11xf32_9_6),
        .p___constant_11x11xf32_9_7(p___constant_11x11xf32_9_7),
        .p___constant_11x11xf32_9_8(p___constant_11x11xf32_9_8),
        .p___constant_11x11xf32_9_9(p___constant_11x11xf32_9_9),
        .p___constant_11xf32_0(p___constant_11xf32_0),
        .p___constant_11xf32_1(p___constant_11xf32_1),
        .p___constant_11xf32_10(p___constant_11xf32_10),
        .p___constant_11xf32_2(p___constant_11xf32_2),
        .p___constant_11xf32_3(p___constant_11xf32_3),
        .p___constant_11xf32_4(p___constant_11xf32_4),
        .p___constant_11xf32_5(p___constant_11xf32_5),
        .p___constant_11xf32_6(p___constant_11xf32_6),
        .p___constant_11xf32_7(p___constant_11xf32_7),
        .p___constant_11xf32_8(p___constant_11xf32_8),
        .p___constant_11xf32_9(p___constant_11xf32_9),
        .output_p_val_313(output_p_val_313)
);


    // Clock generation
initial begin
    forever begin
        #10; // Delay for half a clock cycle (1ns)
        clk <= 1'b0;
        #10; // Delay for half a clock cycle (1ns)
        clk <= 1'b1;
    end
end

    // Initial stimulus
    initial begin
    
    rst = 1;

    p__arg0_0_0 = 12'h6F0;
	p__arg0_0_1 = 12'h6F0;
	p__arg0_0_2 = 12'h6F0;
	p__arg0_0_3 = 12'h6F0;
	p__arg0_0_4 = 12'h6F0;
	p__arg0_0_5 = 12'h6F0;
	p__arg0_0_6 = 12'h6F0;
	p__arg0_0_7 = 12'h6F0;
	p__arg0_0_8 = 12'h6F0;
	p__arg0_0_9 = 12'h6F0;
    p__arg0_0_10 = 12'h6F0;
    p___constant_11x11xf32_0_0 = 12'h6F0;
	p___constant_11x11xf32_0_1 = 12'h6F0;
	p___constant_11x11xf32_0_10 = 12'h6F0;
	p___constant_11x11xf32_0_2 = 12'h6F0;
	p___constant_11x11xf32_0_3 = 12'h6F0;
	p___constant_11x11xf32_0_4 = 12'h6F0;
	p___constant_11x11xf32_0_5 = 12'h6F0;
	p___constant_11x11xf32_0_6 = 12'h6F0;
	p___constant_11x11xf32_0_7 = 12'h6F0;
	p___constant_11x11xf32_0_8 = 12'h6F0;
	p___constant_11x11xf32_0_9 = 12'h6F0;
	p___constant_11x11xf32_10_0 = 12'h6F0;
	p___constant_11x11xf32_10_1 = 12'h6F0;
	p___constant_11x11xf32_10_10 = 12'h6F0;
	p___constant_11x11xf32_10_2 = 12'h6F0;
	p___constant_11x11xf32_10_3 = 12'h6F0;
	p___constant_11x11xf32_10_4 = 12'h6F0;
	p___constant_11x11xf32_10_5 = 12'h6F0;
	p___constant_11x11xf32_10_6 = 12'h6F0;
	p___constant_11x11xf32_10_7 = 12'h6F0;
	p___constant_11x11xf32_10_8 = 12'h6F0;
	p___constant_11x11xf32_10_9 = 12'h6F0;
	p___constant_11x11xf32_1_0 = 12'h6F0;
	p___constant_11x11xf32_1_1 = 12'h6F0;
	p___constant_11x11xf32_1_10 = 12'h6F0;
	p___constant_11x11xf32_1_2 = 12'h6F0;
	p___constant_11x11xf32_1_3 = 12'h6F0;
	p___constant_11x11xf32_1_4 = 12'h6F0;
	p___constant_11x11xf32_1_5 = 12'h6F0;
	p___constant_11x11xf32_1_6 = 12'h6F0;
	p___constant_11x11xf32_1_7 = 12'h6F0;
	p___constant_11x11xf32_1_8 = 12'h6F0;
	p___constant_11x11xf32_1_9 = 12'h6F0;
	p___constant_11x11xf32_2_0 = 12'h6F0;
	p___constant_11x11xf32_2_1 = 12'h6F0;
	p___constant_11x11xf32_2_10 = 12'h6F0;
	p___constant_11x11xf32_2_2 = 12'h6F0;
	p___constant_11x11xf32_2_3 = 12'h6F0;
	p___constant_11x11xf32_2_4 = 12'h6F0;
	p___constant_11x11xf32_2_5 = 12'h6F0;
	p___constant_11x11xf32_2_6 = 12'h6F0;
	p___constant_11x11xf32_2_7 = 12'h6F0;
	p___constant_11x11xf32_2_8 = 12'h6F0;
	p___constant_11x11xf32_2_9 = 12'h6F0;
	p___constant_11x11xf32_3_0 = 12'h6F0;
	p___constant_11x11xf32_3_1 = 12'h6F0;
	p___constant_11x11xf32_3_10 = 12'h6F0;
	p___constant_11x11xf32_3_2 = 12'h6F0;
	p___constant_11x11xf32_3_3 = 12'h6F0;
	p___constant_11x11xf32_3_4 = 12'h6F0;
	p___constant_11x11xf32_3_5 = 12'h6F0;
	p___constant_11x11xf32_3_6 = 12'h6F0;
	p___constant_11x11xf32_3_7 = 12'h6F0;
	p___constant_11x11xf32_3_8 = 12'h6F0;
	p___constant_11x11xf32_3_9 = 12'h6F0;
	p___constant_11x11xf32_4_0 = 12'h6F0;
	p___constant_11x11xf32_4_1 = 12'h6F0;
	p___constant_11x11xf32_4_10 = 12'h6F0;
	p___constant_11x11xf32_4_2 = 12'h6F0;
	p___constant_11x11xf32_4_3 = 12'h6F0;
	p___constant_11x11xf32_4_4 = 12'h6F0;
	p___constant_11x11xf32_4_5 = 12'h6F0;
	p___constant_11x11xf32_4_6 = 12'h6F0;
	p___constant_11x11xf32_4_7 = 12'h6F0;
	p___constant_11x11xf32_4_8 = 12'h6F0;
	p___constant_11x11xf32_4_9 = 12'h6F0;
	p___constant_11x11xf32_5_0 = 12'h6F0;
	p___constant_11x11xf32_5_1 = 12'h6F0;
	p___constant_11x11xf32_5_10 = 12'h6F0;
	p___constant_11x11xf32_5_2 = 12'h6F0;
	p___constant_11x11xf32_5_3 = 12'h6F0;
	p___constant_11x11xf32_5_4 = 12'h6F0;
	p___constant_11x11xf32_5_5 = 12'h6F0;
	p___constant_11x11xf32_5_6 = 12'h6F0;
	p___constant_11x11xf32_5_7 = 12'h6F0;
	p___constant_11x11xf32_5_8 = 12'h6F0;
	p___constant_11x11xf32_5_9 = 12'h6F0;
	p___constant_11x11xf32_6_0 = 12'h6F0;
	p___constant_11x11xf32_6_1 = 12'h6F0;
	p___constant_11x11xf32_6_10 = 12'h6F0;
	p___constant_11x11xf32_6_2 = 12'h6F0;
	p___constant_11x11xf32_6_3 = 12'h6F0;
	p___constant_11x11xf32_6_4 = 12'h6F0;
	p___constant_11x11xf32_6_5 = 12'h6F0;
	p___constant_11x11xf32_6_6 = 12'h6F0;
	p___constant_11x11xf32_6_7 = 12'h6F0;
	p___constant_11x11xf32_6_8 = 12'h6F0;
	p___constant_11x11xf32_6_9 = 12'h6F0;
	p___constant_11x11xf32_7_0 = 12'h6F0;
	p___constant_11x11xf32_7_1 = 12'h6F0;
	p___constant_11x11xf32_7_10 = 12'h6F0;
	p___constant_11x11xf32_7_2 = 12'h6F0;
	p___constant_11x11xf32_7_3 = 12'h6F0;
	p___constant_11x11xf32_7_4 = 12'h6F0;
	p___constant_11x11xf32_7_5 = 12'h6F0;
	p___constant_11x11xf32_7_6 = 12'h6F0;
	p___constant_11x11xf32_7_7 = 12'h6F0;
	p___constant_11x11xf32_7_8 = 12'h6F0;
	p___constant_11x11xf32_7_9 = 12'h6F0;
	p___constant_11x11xf32_8_0 = 12'h6F0;
	p___constant_11x11xf32_8_1 = 12'h6F0;
	p___constant_11x11xf32_8_10 = 12'h6F0;
	p___constant_11x11xf32_8_2 = 12'h6F0;
	p___constant_11x11xf32_8_3 = 12'h6F0;
	p___constant_11x11xf32_8_4 = 12'h6F0;
	p___constant_11x11xf32_8_5 = 12'h6F0;
	p___constant_11x11xf32_8_6 = 12'h6F0;
	p___constant_11x11xf32_8_7 = 12'h6F0;
	p___constant_11x11xf32_8_8 = 12'h6F0;
	p___constant_11x11xf32_8_9 = 12'h6F0;
	p___constant_11x11xf32_9_0 = 12'h6F0;
	p___constant_11x11xf32_9_1 = 12'h6F0;
	p___constant_11x11xf32_9_10 = 12'h6F0;
	p___constant_11x11xf32_9_2 = 12'h6F0;
	p___constant_11x11xf32_9_3 = 12'h6F0;
	p___constant_11x11xf32_9_4 = 12'h6F0;
	p___constant_11x11xf32_9_5 = 12'h6F0;
	p___constant_11x11xf32_9_6 = 12'h6F0;
	p___constant_11x11xf32_9_7 = 12'h6F0;
	p___constant_11x11xf32_9_8 = 12'h6F0;
	p___constant_11x11xf32_9_9 = 12'h6F0;
	p___constant_11xf32_0 = 12'h600;
	p___constant_11xf32_1 = 12'h600;
	p___constant_11xf32_10 = 12'h600;
	p___constant_11xf32_2 = 12'h600;
	p___constant_11xf32_3 = 12'h600;
	p___constant_11xf32_4 = 12'h600;
	p___constant_11xf32_5 = 12'h600;
	p___constant_11xf32_6 = 12'h600;
	p___constant_11xf32_7 = 12'h600;
	p___constant_11xf32_8 = 12'h600;
	p___constant_11xf32_9 = 12'h600;


    #100;

        // Deassert reset
     rst = 0;

        // Add stimulus here if needed

	#5000;

	$display("Output value: %h", output_p_val_313);
	
    end


	

    // Monitor the outputs

endmodule


