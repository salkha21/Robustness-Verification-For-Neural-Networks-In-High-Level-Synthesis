`default_nettype none
module linear (
	clk,
	rst,
	p__arg0_0_0,
	p__arg0_0_1,
	p__arg0_0_10,
	p__arg0_0_2,
	p__arg0_0_3,
	p__arg0_0_4,
	p__arg0_0_5,
	p__arg0_0_6,
	p__arg0_0_7,
	p__arg0_0_8,
	p__arg0_0_9,
	p___constant_11x11xf32_0_0,
	p___constant_11x11xf32_0_1,
	p___constant_11x11xf32_0_10,
	p___constant_11x11xf32_0_2,
	p___constant_11x11xf32_0_3,
	p___constant_11x11xf32_0_4,
	p___constant_11x11xf32_0_5,
	p___constant_11x11xf32_0_6,
	p___constant_11x11xf32_0_7,
	p___constant_11x11xf32_0_8,
	p___constant_11x11xf32_0_9,
	p___constant_11x11xf32_10_0,
	p___constant_11x11xf32_10_1,
	p___constant_11x11xf32_10_10,
	p___constant_11x11xf32_10_2,
	p___constant_11x11xf32_10_3,
	p___constant_11x11xf32_10_4,
	p___constant_11x11xf32_10_5,
	p___constant_11x11xf32_10_6,
	p___constant_11x11xf32_10_7,
	p___constant_11x11xf32_10_8,
	p___constant_11x11xf32_10_9,
	p___constant_11x11xf32_1_0,
	p___constant_11x11xf32_1_1,
	p___constant_11x11xf32_1_10,
	p___constant_11x11xf32_1_2,
	p___constant_11x11xf32_1_3,
	p___constant_11x11xf32_1_4,
	p___constant_11x11xf32_1_5,
	p___constant_11x11xf32_1_6,
	p___constant_11x11xf32_1_7,
	p___constant_11x11xf32_1_8,
	p___constant_11x11xf32_1_9,
	p___constant_11x11xf32_2_0,
	p___constant_11x11xf32_2_1,
	p___constant_11x11xf32_2_10,
	p___constant_11x11xf32_2_2,
	p___constant_11x11xf32_2_3,
	p___constant_11x11xf32_2_4,
	p___constant_11x11xf32_2_5,
	p___constant_11x11xf32_2_6,
	p___constant_11x11xf32_2_7,
	p___constant_11x11xf32_2_8,
	p___constant_11x11xf32_2_9,
	p___constant_11x11xf32_3_0,
	p___constant_11x11xf32_3_1,
	p___constant_11x11xf32_3_10,
	p___constant_11x11xf32_3_2,
	p___constant_11x11xf32_3_3,
	p___constant_11x11xf32_3_4,
	p___constant_11x11xf32_3_5,
	p___constant_11x11xf32_3_6,
	p___constant_11x11xf32_3_7,
	p___constant_11x11xf32_3_8,
	p___constant_11x11xf32_3_9,
	p___constant_11x11xf32_4_0,
	p___constant_11x11xf32_4_1,
	p___constant_11x11xf32_4_10,
	p___constant_11x11xf32_4_2,
	p___constant_11x11xf32_4_3,
	p___constant_11x11xf32_4_4,
	p___constant_11x11xf32_4_5,
	p___constant_11x11xf32_4_6,
	p___constant_11x11xf32_4_7,
	p___constant_11x11xf32_4_8,
	p___constant_11x11xf32_4_9,
	p___constant_11x11xf32_5_0,
	p___constant_11x11xf32_5_1,
	p___constant_11x11xf32_5_10,
	p___constant_11x11xf32_5_2,
	p___constant_11x11xf32_5_3,
	p___constant_11x11xf32_5_4,
	p___constant_11x11xf32_5_5,
	p___constant_11x11xf32_5_6,
	p___constant_11x11xf32_5_7,
	p___constant_11x11xf32_5_8,
	p___constant_11x11xf32_5_9,
	p___constant_11x11xf32_6_0,
	p___constant_11x11xf32_6_1,
	p___constant_11x11xf32_6_10,
	p___constant_11x11xf32_6_2,
	p___constant_11x11xf32_6_3,
	p___constant_11x11xf32_6_4,
	p___constant_11x11xf32_6_5,
	p___constant_11x11xf32_6_6,
	p___constant_11x11xf32_6_7,
	p___constant_11x11xf32_6_8,
	p___constant_11x11xf32_6_9,
	p___constant_11x11xf32_7_0,
	p___constant_11x11xf32_7_1,
	p___constant_11x11xf32_7_10,
	p___constant_11x11xf32_7_2,
	p___constant_11x11xf32_7_3,
	p___constant_11x11xf32_7_4,
	p___constant_11x11xf32_7_5,
	p___constant_11x11xf32_7_6,
	p___constant_11x11xf32_7_7,
	p___constant_11x11xf32_7_8,
	p___constant_11x11xf32_7_9,
	p___constant_11x11xf32_8_0,
	p___constant_11x11xf32_8_1,
	p___constant_11x11xf32_8_10,
	p___constant_11x11xf32_8_2,
	p___constant_11x11xf32_8_3,
	p___constant_11x11xf32_8_4,
	p___constant_11x11xf32_8_5,
	p___constant_11x11xf32_8_6,
	p___constant_11x11xf32_8_7,
	p___constant_11x11xf32_8_8,
	p___constant_11x11xf32_8_9,
	p___constant_11x11xf32_9_0,
	p___constant_11x11xf32_9_1,
	p___constant_11x11xf32_9_10,
	p___constant_11x11xf32_9_2,
	p___constant_11x11xf32_9_3,
	p___constant_11x11xf32_9_4,
	p___constant_11x11xf32_9_5,
	p___constant_11x11xf32_9_6,
	p___constant_11x11xf32_9_7,
	p___constant_11x11xf32_9_8,
	p___constant_11x11xf32_9_9,
	p___constant_11xf32_0,
	p___constant_11xf32_1,
	p___constant_11xf32_10,
	p___constant_11xf32_2,
	p___constant_11xf32_3,
	p___constant_11xf32_4,
	p___constant_11xf32_5,
	p___constant_11xf32_6,
	p___constant_11xf32_7,
	p___constant_11xf32_8,
	p___constant_11xf32_9,
	output_p_val_313
);
	input wire clk;
	input wire rst;
	input wire [11:0] p__arg0_0_0;
	input wire [11:0] p__arg0_0_1;
	input wire [11:0] p__arg0_0_10;
	input wire [11:0] p__arg0_0_2;
	input wire [11:0] p__arg0_0_3;
	input wire [11:0] p__arg0_0_4;
	input wire [11:0] p__arg0_0_5;
	input wire [11:0] p__arg0_0_6;
	input wire [11:0] p__arg0_0_7;
	input wire [11:0] p__arg0_0_8;
	input wire [11:0] p__arg0_0_9;
	input wire [11:0] p___constant_11x11xf32_0_0;
	input wire [11:0] p___constant_11x11xf32_0_1;
	input wire [11:0] p___constant_11x11xf32_0_10;
	input wire [11:0] p___constant_11x11xf32_0_2;
	input wire [11:0] p___constant_11x11xf32_0_3;
	input wire [11:0] p___constant_11x11xf32_0_4;
	input wire [11:0] p___constant_11x11xf32_0_5;
	input wire [11:0] p___constant_11x11xf32_0_6;
	input wire [11:0] p___constant_11x11xf32_0_7;
	input wire [11:0] p___constant_11x11xf32_0_8;
	input wire [11:0] p___constant_11x11xf32_0_9;
	input wire [11:0] p___constant_11x11xf32_10_0;
	input wire [11:0] p___constant_11x11xf32_10_1;
	input wire [11:0] p___constant_11x11xf32_10_10;
	input wire [11:0] p___constant_11x11xf32_10_2;
	input wire [11:0] p___constant_11x11xf32_10_3;
	input wire [11:0] p___constant_11x11xf32_10_4;
	input wire [11:0] p___constant_11x11xf32_10_5;
	input wire [11:0] p___constant_11x11xf32_10_6;
	input wire [11:0] p___constant_11x11xf32_10_7;
	input wire [11:0] p___constant_11x11xf32_10_8;
	input wire [11:0] p___constant_11x11xf32_10_9;
	input wire [11:0] p___constant_11x11xf32_1_0;
	input wire [11:0] p___constant_11x11xf32_1_1;
	input wire [11:0] p___constant_11x11xf32_1_10;
	input wire [11:0] p___constant_11x11xf32_1_2;
	input wire [11:0] p___constant_11x11xf32_1_3;
	input wire [11:0] p___constant_11x11xf32_1_4;
	input wire [11:0] p___constant_11x11xf32_1_5;
	input wire [11:0] p___constant_11x11xf32_1_6;
	input wire [11:0] p___constant_11x11xf32_1_7;
	input wire [11:0] p___constant_11x11xf32_1_8;
	input wire [11:0] p___constant_11x11xf32_1_9;
	input wire [11:0] p___constant_11x11xf32_2_0;
	input wire [11:0] p___constant_11x11xf32_2_1;
	input wire [11:0] p___constant_11x11xf32_2_10;
	input wire [11:0] p___constant_11x11xf32_2_2;
	input wire [11:0] p___constant_11x11xf32_2_3;
	input wire [11:0] p___constant_11x11xf32_2_4;
	input wire [11:0] p___constant_11x11xf32_2_5;
	input wire [11:0] p___constant_11x11xf32_2_6;
	input wire [11:0] p___constant_11x11xf32_2_7;
	input wire [11:0] p___constant_11x11xf32_2_8;
	input wire [11:0] p___constant_11x11xf32_2_9;
	input wire [11:0] p___constant_11x11xf32_3_0;
	input wire [11:0] p___constant_11x11xf32_3_1;
	input wire [11:0] p___constant_11x11xf32_3_10;
	input wire [11:0] p___constant_11x11xf32_3_2;
	input wire [11:0] p___constant_11x11xf32_3_3;
	input wire [11:0] p___constant_11x11xf32_3_4;
	input wire [11:0] p___constant_11x11xf32_3_5;
	input wire [11:0] p___constant_11x11xf32_3_6;
	input wire [11:0] p___constant_11x11xf32_3_7;
	input wire [11:0] p___constant_11x11xf32_3_8;
	input wire [11:0] p___constant_11x11xf32_3_9;
	input wire [11:0] p___constant_11x11xf32_4_0;
	input wire [11:0] p___constant_11x11xf32_4_1;
	input wire [11:0] p___constant_11x11xf32_4_10;
	input wire [11:0] p___constant_11x11xf32_4_2;
	input wire [11:0] p___constant_11x11xf32_4_3;
	input wire [11:0] p___constant_11x11xf32_4_4;
	input wire [11:0] p___constant_11x11xf32_4_5;
	input wire [11:0] p___constant_11x11xf32_4_6;
	input wire [11:0] p___constant_11x11xf32_4_7;
	input wire [11:0] p___constant_11x11xf32_4_8;
	input wire [11:0] p___constant_11x11xf32_4_9;
	input wire [11:0] p___constant_11x11xf32_5_0;
	input wire [11:0] p___constant_11x11xf32_5_1;
	input wire [11:0] p___constant_11x11xf32_5_10;
	input wire [11:0] p___constant_11x11xf32_5_2;
	input wire [11:0] p___constant_11x11xf32_5_3;
	input wire [11:0] p___constant_11x11xf32_5_4;
	input wire [11:0] p___constant_11x11xf32_5_5;
	input wire [11:0] p___constant_11x11xf32_5_6;
	input wire [11:0] p___constant_11x11xf32_5_7;
	input wire [11:0] p___constant_11x11xf32_5_8;
	input wire [11:0] p___constant_11x11xf32_5_9;
	input wire [11:0] p___constant_11x11xf32_6_0;
	input wire [11:0] p___constant_11x11xf32_6_1;
	input wire [11:0] p___constant_11x11xf32_6_10;
	input wire [11:0] p___constant_11x11xf32_6_2;
	input wire [11:0] p___constant_11x11xf32_6_3;
	input wire [11:0] p___constant_11x11xf32_6_4;
	input wire [11:0] p___constant_11x11xf32_6_5;
	input wire [11:0] p___constant_11x11xf32_6_6;
	input wire [11:0] p___constant_11x11xf32_6_7;
	input wire [11:0] p___constant_11x11xf32_6_8;
	input wire [11:0] p___constant_11x11xf32_6_9;
	input wire [11:0] p___constant_11x11xf32_7_0;
	input wire [11:0] p___constant_11x11xf32_7_1;
	input wire [11:0] p___constant_11x11xf32_7_10;
	input wire [11:0] p___constant_11x11xf32_7_2;
	input wire [11:0] p___constant_11x11xf32_7_3;
	input wire [11:0] p___constant_11x11xf32_7_4;
	input wire [11:0] p___constant_11x11xf32_7_5;
	input wire [11:0] p___constant_11x11xf32_7_6;
	input wire [11:0] p___constant_11x11xf32_7_7;
	input wire [11:0] p___constant_11x11xf32_7_8;
	input wire [11:0] p___constant_11x11xf32_7_9;
	input wire [11:0] p___constant_11x11xf32_8_0;
	input wire [11:0] p___constant_11x11xf32_8_1;
	input wire [11:0] p___constant_11x11xf32_8_10;
	input wire [11:0] p___constant_11x11xf32_8_2;
	input wire [11:0] p___constant_11x11xf32_8_3;
	input wire [11:0] p___constant_11x11xf32_8_4;
	input wire [11:0] p___constant_11x11xf32_8_5;
	input wire [11:0] p___constant_11x11xf32_8_6;
	input wire [11:0] p___constant_11x11xf32_8_7;
	input wire [11:0] p___constant_11x11xf32_8_8;
	input wire [11:0] p___constant_11x11xf32_8_9;
	input wire [11:0] p___constant_11x11xf32_9_0;
	input wire [11:0] p___constant_11x11xf32_9_1;
	input wire [11:0] p___constant_11x11xf32_9_10;
	input wire [11:0] p___constant_11x11xf32_9_2;
	input wire [11:0] p___constant_11x11xf32_9_3;
	input wire [11:0] p___constant_11x11xf32_9_4;
	input wire [11:0] p___constant_11x11xf32_9_5;
	input wire [11:0] p___constant_11x11xf32_9_6;
	input wire [11:0] p___constant_11x11xf32_9_7;
	input wire [11:0] p___constant_11x11xf32_9_8;
	input wire [11:0] p___constant_11x11xf32_9_9;
	input wire [11:0] p___constant_11xf32_0;
	input wire [11:0] p___constant_11xf32_1;
	input wire [11:0] p___constant_11xf32_10;
	input wire [11:0] p___constant_11xf32_2;
	input wire [11:0] p___constant_11xf32_3;
	input wire [11:0] p___constant_11xf32_4;
	input wire [11:0] p___constant_11xf32_5;
	input wire [11:0] p___constant_11xf32_6;
	input wire [11:0] p___constant_11xf32_7;
	input wire [11:0] p___constant_11xf32_8;
	input wire [11:0] p___constant_11xf32_9;
	output wire [11:0] output_p_val_313;



reg [11:0] p_val_106;

reg [11:0] p_val_107;

reg [11:0] p_val_130;

reg [11:0] p_val_131;

reg [11:0] p_val_154;

reg [11:0] p_val_155;

reg [11:0] p_val_178;

reg [11:0] p_val_179;

reg [11:0] p_val_202;

reg [11:0] p_val_203;

reg [11:0] p_val_226;

reg [11:0] p_val_227;

reg [11:0] p_val_250;

reg [11:0] p_val_251;

reg [11:0] p_val_274;

reg [11:0] p_val_275;

reg [11:0] p_val_276;

reg [11:0] p_val_277;

reg [11:0] p_val_278;

reg [11:0] p_val_279;

reg [11:0] p_val_280;

reg [11:0] p_val_281;

reg [11:0] p_val_282;

reg [11:0] p_val_283;

reg [11:0] p_val_284;

reg [11:0] p_val_285;

reg [11:0] p_val_286;

reg [11:0] p_val_287;

reg [11:0] p_val_288;

reg [11:0] p_val_289;

reg [11:0] p_val_290;

reg [11:0] p_val_291;

reg [11:0] p_val_292;

reg [11:0] p_val_293;

reg [11:0] p_val_294;

reg [11:0] p_val_295;

reg [11:0] p_val_296;

reg [11:0] p_val_297;

reg [11:0] p_val_299;

reg [11:0] p_val_300;

reg [11:0] p_val_301;

reg [11:0] p_val_302;

reg [11:0] p_val_303;

reg [11:0] p_val_304;

reg [11:0] p_val_305;

reg [11:0] p_val_306;

reg [11:0] p_val_307;

reg [11:0] p_val_308;

reg [11:0] p_val_309;

reg [11:0] p_val_310;

reg [11:0] p_val_311;

reg [11:0] p_val_312;

reg [11:0] p_val_313;

reg [11:0] p_val_34;

reg [11:0] p_val_35;

reg [11:0] p_val_58;

reg [11:0] p_val_59;

reg [11:0] p_val_82;

reg [11:0] p_val_83;

reg [11:0] p_val_cst_0_point_0000000000000000000000000 = 12'b000000000000; // 0.0

parameter fsm_state01 = 56'd1;
parameter fsm_state02 = 56'd2;
parameter fsm_state03 = 56'd4;
parameter fsm_state04 = 56'd8;
parameter fsm_state05 = 56'd16;
parameter fsm_state06 = 56'd32;
parameter fsm_state07 = 56'd64;
parameter fsm_state08 = 56'd128;
parameter fsm_state09 = 56'd256;
parameter fsm_state10 = 56'd512;
parameter fsm_state11 = 56'd1024;
parameter fsm_state12 = 56'd2048;
parameter fsm_state13 = 56'd4096;
parameter fsm_state14 = 56'd8192;
parameter fsm_state15 = 56'd16384;
parameter fsm_state16 = 56'd32768;
parameter fsm_state17 = 56'd65536;
parameter fsm_state18 = 56'd131072;
parameter fsm_state19 = 56'd262144;
parameter fsm_state20 = 56'd524288;
parameter fsm_state21 = 56'd1048576;
parameter fsm_state22 = 56'd2097152;
parameter fsm_state23 = 56'd4194304;
parameter fsm_state24 = 56'd8388608;
parameter fsm_state25 = 56'd16777216;
parameter fsm_state26 = 56'd33554432;
parameter fsm_state27 = 56'd67108864;
parameter fsm_state28 = 56'd134217728;
parameter fsm_state29 = 56'd268435456;
parameter fsm_state30 = 56'd536870912;
parameter fsm_state31 = 56'd1073741824;
parameter fsm_state32 = 56'd2147483648;
parameter fsm_state33 = 56'd4294967296;
parameter fsm_state34 = 56'd8589934592;
parameter fsm_state35 = 56'd17179869184;
parameter fsm_state36 = 56'd34359738368;
parameter fsm_state37 = 56'd68719476736;
parameter fsm_state38 = 56'd137438953472;
parameter fsm_state39 = 56'd274877906944;
parameter fsm_state40 = 56'd549755813888;
parameter fsm_state41 = 56'd1099511627776;
parameter fsm_state42 = 56'd2199023255552;
parameter fsm_state43 = 56'd4398046511104;
parameter fsm_state44 = 56'd8796093022208;
parameter fsm_state45 = 56'd17592186044416;
parameter fsm_state46 = 56'd35184372088832;
parameter fsm_state47 = 56'd70368744177664;
parameter fsm_state48 = 56'd140737488355328;
parameter fsm_state49 = 56'd281474976710656;
parameter fsm_state50 = 56'd562949953421312;
parameter fsm_state51 = 56'd1125899906842624;
parameter fsm_state52 = 56'd2251799813685248;
parameter fsm_state53 = 56'd4503599627370496;
parameter fsm_state54 = 56'd9007199254740992;
parameter fsm_state55 = 56'd18014398509481984;

(* max_fanout = 50, fsm_encoding = "none" *) reg [55:0] current_fsm;
reg [55:0] next_state_fsm;

wire current_fsm_state01;
wire current_fsm_state02;
wire current_fsm_state03;
wire current_fsm_state04;
wire current_fsm_state05;
wire current_fsm_state06;
wire current_fsm_state07;
wire current_fsm_state08;
wire current_fsm_state09;
wire current_fsm_state10;
wire current_fsm_state11;
wire current_fsm_state12;
wire current_fsm_state13;
wire current_fsm_state14;
wire current_fsm_state15;
wire current_fsm_state16;
wire current_fsm_state17;
wire current_fsm_state18;
wire current_fsm_state19;
wire current_fsm_state20;
wire current_fsm_state21;
wire current_fsm_state22;
wire current_fsm_state23;
wire current_fsm_state24;
wire current_fsm_state25;
wire current_fsm_state26;
wire current_fsm_state27;
wire current_fsm_state28;
wire current_fsm_state29;
wire current_fsm_state30;
wire current_fsm_state31;
wire current_fsm_state32;
wire current_fsm_state33;
wire current_fsm_state34;
wire current_fsm_state35;
wire current_fsm_state36;
wire current_fsm_state37;
wire current_fsm_state38;
wire current_fsm_state39;
wire current_fsm_state40;
wire current_fsm_state41;
wire current_fsm_state42;
wire current_fsm_state43;
wire current_fsm_state44;
wire current_fsm_state45;
wire current_fsm_state46;
wire current_fsm_state47;
wire current_fsm_state48;
wire current_fsm_state49;
wire current_fsm_state50;
wire current_fsm_state51;
wire current_fsm_state52;
wire current_fsm_state53;
wire current_fsm_state54;
wire current_fsm_state55;

reg [11:0] fadd_0_0_0_0_0_x;
reg [11:0] fadd_0_0_0_0_0_y;
wire [11:0] fadd_0_0_0_0_0_r;
fadd #(1) fadd_0_0_0_0_0(
    .clk(clk),
    .X(fadd_0_0_0_0_0_x),
    .Y(fadd_0_0_0_0_0_y),
    .R(fadd_0_0_0_0_0_r)
);


reg [11:0] fmul_0_0_0_0_0_x;
reg [11:0] fmul_0_0_0_0_0_y;
wire [11:0] fmul_0_0_0_0_0_r;
fmul #(1) fmul_0_0_0_0_0(
    .clk(clk),
    .X(fmul_0_0_0_0_0_x),
    .Y(fmul_0_0_0_0_0_y),
    .R(fmul_0_0_0_0_0_r)
);


reg [11:0] fadd_0_0_0_0_1_x;
reg [11:0] fadd_0_0_0_0_1_y;
wire [11:0] fadd_0_0_0_0_1_r;
fadd #(1) fadd_0_0_0_0_1(
    .clk(clk),
    .X(fadd_0_0_0_0_1_x),
    .Y(fadd_0_0_0_0_1_y),
    .R(fadd_0_0_0_0_1_r)
);


reg [11:0] fmul_0_0_0_0_1_x;
reg [11:0] fmul_0_0_0_0_1_y;
wire [11:0] fmul_0_0_0_0_1_r;
fmul #(1) fmul_0_0_0_0_1(
    .clk(clk),
    .X(fmul_0_0_0_0_1_x),
    .Y(fmul_0_0_0_0_1_y),
    .R(fmul_0_0_0_0_1_r)
);


reg [11:0] fadd_0_0_0_0_2_x;
reg [11:0] fadd_0_0_0_0_2_y;
wire [11:0] fadd_0_0_0_0_2_r;
fadd #(1) fadd_0_0_0_0_2(
    .clk(clk),
    .X(fadd_0_0_0_0_2_x),
    .Y(fadd_0_0_0_0_2_y),
    .R(fadd_0_0_0_0_2_r)
);


reg [11:0] fmul_0_0_0_0_2_x;
reg [11:0] fmul_0_0_0_0_2_y;
wire [11:0] fmul_0_0_0_0_2_r;
fmul #(1) fmul_0_0_0_0_2(
    .clk(clk),
    .X(fmul_0_0_0_0_2_x),
    .Y(fmul_0_0_0_0_2_y),
    .R(fmul_0_0_0_0_2_r)
);


reg [11:0] fadd_0_0_0_0_3_x;
reg [11:0] fadd_0_0_0_0_3_y;
wire [11:0] fadd_0_0_0_0_3_r;
fadd #(1) fadd_0_0_0_0_3(
    .clk(clk),
    .X(fadd_0_0_0_0_3_x),
    .Y(fadd_0_0_0_0_3_y),
    .R(fadd_0_0_0_0_3_r)
);


reg [11:0] fmul_0_0_0_0_3_x;
reg [11:0] fmul_0_0_0_0_3_y;
wire [11:0] fmul_0_0_0_0_3_r;
fmul #(1) fmul_0_0_0_0_3(
    .clk(clk),
    .X(fmul_0_0_0_0_3_x),
    .Y(fmul_0_0_0_0_3_y),
    .R(fmul_0_0_0_0_3_r)
);


reg [11:0] fadd_0_0_0_0_4_x;
reg [11:0] fadd_0_0_0_0_4_y;
wire [11:0] fadd_0_0_0_0_4_r;
fadd #(1) fadd_0_0_0_0_4(
    .clk(clk),
    .X(fadd_0_0_0_0_4_x),
    .Y(fadd_0_0_0_0_4_y),
    .R(fadd_0_0_0_0_4_r)
);


reg [11:0] fmul_0_0_0_0_4_x;
reg [11:0] fmul_0_0_0_0_4_y;
wire [11:0] fmul_0_0_0_0_4_r;
fmul #(1) fmul_0_0_0_0_4(
    .clk(clk),
    .X(fmul_0_0_0_0_4_x),
    .Y(fmul_0_0_0_0_4_y),
    .R(fmul_0_0_0_0_4_r)
);


reg [11:0] fadd_0_0_0_0_5_x;
reg [11:0] fadd_0_0_0_0_5_y;
wire [11:0] fadd_0_0_0_0_5_r;
fadd #(1) fadd_0_0_0_0_5(
    .clk(clk),
    .X(fadd_0_0_0_0_5_x),
    .Y(fadd_0_0_0_0_5_y),
    .R(fadd_0_0_0_0_5_r)
);


reg [11:0] fmul_0_0_0_0_5_x;
reg [11:0] fmul_0_0_0_0_5_y;
wire [11:0] fmul_0_0_0_0_5_r;
fmul #(1) fmul_0_0_0_0_5(
    .clk(clk),
    .X(fmul_0_0_0_0_5_x),
    .Y(fmul_0_0_0_0_5_y),
    .R(fmul_0_0_0_0_5_r)
);


reg [11:0] fadd_0_0_0_0_6_x;
reg [11:0] fadd_0_0_0_0_6_y;
wire [11:0] fadd_0_0_0_0_6_r;
fadd #(1) fadd_0_0_0_0_6(
    .clk(clk),
    .X(fadd_0_0_0_0_6_x),
    .Y(fadd_0_0_0_0_6_y),
    .R(fadd_0_0_0_0_6_r)
);


reg [11:0] fmul_0_0_0_0_6_x;
reg [11:0] fmul_0_0_0_0_6_y;
wire [11:0] fmul_0_0_0_0_6_r;
fmul #(1) fmul_0_0_0_0_6(
    .clk(clk),
    .X(fmul_0_0_0_0_6_x),
    .Y(fmul_0_0_0_0_6_y),
    .R(fmul_0_0_0_0_6_r)
);


reg [11:0] fadd_0_0_0_0_7_x;
reg [11:0] fadd_0_0_0_0_7_y;
wire [11:0] fadd_0_0_0_0_7_r;
fadd #(1) fadd_0_0_0_0_7(
    .clk(clk),
    .X(fadd_0_0_0_0_7_x),
    .Y(fadd_0_0_0_0_7_y),
    .R(fadd_0_0_0_0_7_r)
);


reg [11:0] fmul_0_0_0_0_7_x;
reg [11:0] fmul_0_0_0_0_7_y;
wire [11:0] fmul_0_0_0_0_7_r;
fmul #(1) fmul_0_0_0_0_7(
    .clk(clk),
    .X(fmul_0_0_0_0_7_x),
    .Y(fmul_0_0_0_0_7_y),
    .R(fmul_0_0_0_0_7_r)
);


reg [11:0] fadd_0_0_0_0_8_x;
reg [11:0] fadd_0_0_0_0_8_y;
wire [11:0] fadd_0_0_0_0_8_r;
fadd #(1) fadd_0_0_0_0_8(
    .clk(clk),
    .X(fadd_0_0_0_0_8_x),
    .Y(fadd_0_0_0_0_8_y),
    .R(fadd_0_0_0_0_8_r)
);


reg [11:0] fmul_0_0_0_0_8_x;
reg [11:0] fmul_0_0_0_0_8_y;
wire [11:0] fmul_0_0_0_0_8_r;
fmul #(1) fmul_0_0_0_0_8(
    .clk(clk),
    .X(fmul_0_0_0_0_8_x),
    .Y(fmul_0_0_0_0_8_y),
    .R(fmul_0_0_0_0_8_r)
);


reg [11:0] fadd_0_0_0_0_9_x;
reg [11:0] fadd_0_0_0_0_9_y;
wire [11:0] fadd_0_0_0_0_9_r;
fadd #(1) fadd_0_0_0_0_9(
    .clk(clk),
    .X(fadd_0_0_0_0_9_x),
    .Y(fadd_0_0_0_0_9_y),
    .R(fadd_0_0_0_0_9_r)
);


reg [11:0] fmul_0_0_0_0_9_x;
reg [11:0] fmul_0_0_0_0_9_y;
wire [11:0] fmul_0_0_0_0_9_r;
fmul #(1) fmul_0_0_0_0_9(
    .clk(clk),
    .X(fmul_0_0_0_0_9_x),
    .Y(fmul_0_0_0_0_9_y),
    .R(fmul_0_0_0_0_9_r)
);


reg [11:0] fadd_0_0_0_0_10_x;
reg [11:0] fadd_0_0_0_0_10_y;
wire [11:0] fadd_0_0_0_0_10_r;
fadd #(1) fadd_0_0_0_0_10(
    .clk(clk),
    .X(fadd_0_0_0_0_10_x),
    .Y(fadd_0_0_0_0_10_y),
    .R(fadd_0_0_0_0_10_r)
);


reg [11:0] fmul_0_0_0_0_10_x;
reg [11:0] fmul_0_0_0_0_10_y;
wire [11:0] fmul_0_0_0_0_10_r;
fmul #(1) fmul_0_0_0_0_10(
    .clk(clk),
    .X(fmul_0_0_0_0_10_x),
    .Y(fmul_0_0_0_0_10_y),
    .R(fmul_0_0_0_0_10_r)
);


always @ (posedge clk) begin

	// p_val_34 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_0_0, p__arg0_0_1, p___constant_11x11xf32_0_1, p__arg0_0_2, p___constant_11x11xf32_0_2, p__arg0_0_3, p___constant_11x11xf32_0_3, p__arg0_0_4, p___constant_11x11xf32_0_4, p__arg0_0_5, p___constant_11x11xf32_0_5, p__arg0_0_6, p___constant_11x11xf32_0_6, p__arg0_0_7, p___constant_11x11xf32_0_7, p__arg0_0_8, p___constant_11x11xf32_0_8, p__arg0_0_9, p___constant_11x11xf32_0_9, p__arg0_0_10, p___constant_11x11xf32_0_10) {  pe = "(0, 0, 0, 0, 0)", opr = "fmac", op_id = "1", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 start
	if (1'b1 == current_fsm_state01) begin
	    fmul_0_0_0_0_0_x <= p__arg0_0_0;
	    fmul_0_0_0_0_0_y <= p___constant_11x11xf32_0_0;
	end
	if (1'b1 == current_fsm_state03) begin
	    fadd_0_0_0_0_0_x <= p_val_cst_0_point_0000000000000000000000000;
	    fadd_0_0_0_0_0_y <= fmul_0_0_0_0_0_r;
	end

	if (1'b1 == current_fsm_state04) begin
	    fmul_0_0_0_0_0_x <= p__arg0_0_1;
	    fmul_0_0_0_0_0_y <= p___constant_11x11xf32_0_1;
	end
	if (1'b1 == current_fsm_state06) begin
	    fadd_0_0_0_0_0_x <= fadd_0_0_0_0_0_r;
	    fadd_0_0_0_0_0_y <= fmul_0_0_0_0_0_r;
	end

	if (1'b1 == current_fsm_state07) begin
	    fmul_0_0_0_0_0_x <= p__arg0_0_2;
	    fmul_0_0_0_0_0_y <= p___constant_11x11xf32_0_2;
	end
	if (1'b1 == current_fsm_state09) begin
	    fadd_0_0_0_0_0_x <= fadd_0_0_0_0_0_r;
	    fadd_0_0_0_0_0_y <= fmul_0_0_0_0_0_r;
	end

	if (1'b1 == current_fsm_state10) begin
	    fmul_0_0_0_0_0_x <= p__arg0_0_3;
	    fmul_0_0_0_0_0_y <= p___constant_11x11xf32_0_3;
	end
	if (1'b1 == current_fsm_state12) begin
	    fadd_0_0_0_0_0_x <= fadd_0_0_0_0_0_r;
	    fadd_0_0_0_0_0_y <= fmul_0_0_0_0_0_r;
	end

	if (1'b1 == current_fsm_state13) begin
	    fmul_0_0_0_0_0_x <= p__arg0_0_4;
	    fmul_0_0_0_0_0_y <= p___constant_11x11xf32_0_4;
	end
	if (1'b1 == current_fsm_state15) begin
	    fadd_0_0_0_0_0_x <= fadd_0_0_0_0_0_r;
	    fadd_0_0_0_0_0_y <= fmul_0_0_0_0_0_r;
	end

	if (1'b1 == current_fsm_state16) begin
	    fmul_0_0_0_0_0_x <= p__arg0_0_5;
	    fmul_0_0_0_0_0_y <= p___constant_11x11xf32_0_5;
	end
	if (1'b1 == current_fsm_state18) begin
	    fadd_0_0_0_0_0_x <= fadd_0_0_0_0_0_r;
	    fadd_0_0_0_0_0_y <= fmul_0_0_0_0_0_r;
	end

	if (1'b1 == current_fsm_state19) begin
	    fmul_0_0_0_0_0_x <= p__arg0_0_6;
	    fmul_0_0_0_0_0_y <= p___constant_11x11xf32_0_6;
	end
	if (1'b1 == current_fsm_state21) begin
	    fadd_0_0_0_0_0_x <= fadd_0_0_0_0_0_r;
	    fadd_0_0_0_0_0_y <= fmul_0_0_0_0_0_r;
	end

	if (1'b1 == current_fsm_state22) begin
	    fmul_0_0_0_0_0_x <= p__arg0_0_7;
	    fmul_0_0_0_0_0_y <= p___constant_11x11xf32_0_7;
	end
	if (1'b1 == current_fsm_state24) begin
	    fadd_0_0_0_0_0_x <= fadd_0_0_0_0_0_r;
	    fadd_0_0_0_0_0_y <= fmul_0_0_0_0_0_r;
	end

	if (1'b1 == current_fsm_state25) begin
	    fmul_0_0_0_0_0_x <= p__arg0_0_8;
	    fmul_0_0_0_0_0_y <= p___constant_11x11xf32_0_8;
	end
	if (1'b1 == current_fsm_state27) begin
	    fadd_0_0_0_0_0_x <= fadd_0_0_0_0_0_r;
	    fadd_0_0_0_0_0_y <= fmul_0_0_0_0_0_r;
	end

	if (1'b1 == current_fsm_state28) begin
	    fmul_0_0_0_0_0_x <= p__arg0_0_9;
	    fmul_0_0_0_0_0_y <= p___constant_11x11xf32_0_9;
	end
	if (1'b1 == current_fsm_state30) begin
	    fadd_0_0_0_0_0_x <= fadd_0_0_0_0_0_r;
	    fadd_0_0_0_0_0_y <= fmul_0_0_0_0_0_r;
	end

	if (1'b1 == current_fsm_state31) begin
	    fmul_0_0_0_0_0_x <= p__arg0_0_10;
	    fmul_0_0_0_0_0_y <= p___constant_11x11xf32_0_10;
	end
	if (1'b1 == current_fsm_state33) begin
	    fadd_0_0_0_0_0_x <= fadd_0_0_0_0_0_r;
	    fadd_0_0_0_0_0_y <= fmul_0_0_0_0_0_r;
	end

	// p_val_34 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_0_0, p__arg0_0_1, p___constant_11x11xf32_0_1, p__arg0_0_2, p___constant_11x11xf32_0_2, p__arg0_0_3, p___constant_11x11xf32_0_3, p__arg0_0_4, p___constant_11x11xf32_0_4, p__arg0_0_5, p___constant_11x11xf32_0_5, p__arg0_0_6, p___constant_11x11xf32_0_6, p__arg0_0_7, p___constant_11x11xf32_0_7, p__arg0_0_8, p___constant_11x11xf32_0_8, p__arg0_0_9, p___constant_11x11xf32_0_9, p__arg0_0_10, p___constant_11x11xf32_0_10) {  pe = "(0, 0, 0, 0, 0)", opr = "fmac", op_id = "1", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 end


	// p_val_35 = "copy" (p_val_34) {  pe = "(0, 0, 0, 0, 0)", opr = "copy", op_id = "2", start_time = "36"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state36) begin
	    p_val_35 <= fadd_0_0_0_0_0_r;
	end
	// p_val_35 = "copy" (p_val_34) {  pe = "(0, 0, 0, 0, 0)", opr = "copy", op_id = "2", start_time = "36"  } : (f32) -> f32 end


	// p_val_276 = "fadd" (p_val_35, p___constant_11xf32_0) {  pe = "(0, 0, 0, 0, 0)", opr = "fadd", op_id = "23", start_time = "37"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state37) begin
	    fadd_0_0_0_0_0_x <= p_val_35;
	    fadd_0_0_0_0_0_y <= p___constant_11xf32_0;
	end
	// p_val_276 = "fadd" (p_val_35, p___constant_11xf32_0) {  pe = "(0, 0, 0, 0, 0)", opr = "fadd", op_id = "23", start_time = "37"  } : (f32, f32) -> f32 end


	// p_val_287 = "copy" (p_val_276) {  pe = "(0, 0, 0, 0, 0)", opr = "copy", op_id = "34", start_time = "40"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state40) begin
	    p_val_287 <= fadd_0_0_0_0_0_r;
	end
	// p_val_287 = "copy" (p_val_276) {  pe = "(0, 0, 0, 0, 0)", opr = "copy", op_id = "34", start_time = "40"  } : (f32) -> f32 end


	// p_val_299 = "fadd" (p_val_287, p_val_288) {  pe = "(0, 0, 0, 0, 0)", opr = "fadd", op_id = "45", start_time = "41"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state41) begin
	    fadd_0_0_0_0_0_x <= p_val_287;
	    fadd_0_0_0_0_0_y <= p_val_288;
	end
	// p_val_299 = "fadd" (p_val_287, p_val_288) {  pe = "(0, 0, 0, 0, 0)", opr = "fadd", op_id = "45", start_time = "41"  } : (f32, f32) -> f32 end


	// p_val_303 = "fadd" (p_val_299, p_val_300) {  pe = "(0, 0, 0, 0, 0)", opr = "fadd", op_id = "49", start_time = "44"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state44) begin
	    fadd_0_0_0_0_0_x <= fadd_0_0_0_0_0_r;
	    fadd_0_0_0_0_0_y <= fadd_0_0_0_0_2_r;
	end
	// p_val_303 = "fadd" (p_val_299, p_val_300) {  pe = "(0, 0, 0, 0, 0)", opr = "fadd", op_id = "49", start_time = "44"  } : (f32, f32) -> f32 end


	// p_val_305 = "fadd" (p_val_303, p_val_304) {  pe = "(0, 0, 0, 0, 0)", opr = "fadd", op_id = "51", start_time = "47"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state47) begin
	    fadd_0_0_0_0_0_x <= fadd_0_0_0_0_0_r;
	    fadd_0_0_0_0_0_y <= fadd_0_0_0_0_4_r;
	end
	// p_val_305 = "fadd" (p_val_303, p_val_304) {  pe = "(0, 0, 0, 0, 0)", opr = "fadd", op_id = "51", start_time = "47"  } : (f32, f32) -> f32 end

end

always @ (posedge clk) begin

	// p_val_58 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_1_0, p__arg0_0_1, p___constant_11x11xf32_1_1, p__arg0_0_2, p___constant_11x11xf32_1_2, p__arg0_0_3, p___constant_11x11xf32_1_3, p__arg0_0_4, p___constant_11x11xf32_1_4, p__arg0_0_5, p___constant_11x11xf32_1_5, p__arg0_0_6, p___constant_11x11xf32_1_6, p__arg0_0_7, p___constant_11x11xf32_1_7, p__arg0_0_8, p___constant_11x11xf32_1_8, p__arg0_0_9, p___constant_11x11xf32_1_9, p__arg0_0_10, p___constant_11x11xf32_1_10) {  pe = "(0, 0, 0, 0, 1)", opr = "fmac", op_id = "3", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 start
	if (1'b1 == current_fsm_state01) begin
	    fmul_0_0_0_0_1_x <= p__arg0_0_0;
	    fmul_0_0_0_0_1_y <= p___constant_11x11xf32_1_0;
	end
	if (1'b1 == current_fsm_state03) begin
	    fadd_0_0_0_0_1_x <= p_val_cst_0_point_0000000000000000000000000;
	    fadd_0_0_0_0_1_y <= fmul_0_0_0_0_1_r;
	end

	if (1'b1 == current_fsm_state04) begin
	    fmul_0_0_0_0_1_x <= p__arg0_0_1;
	    fmul_0_0_0_0_1_y <= p___constant_11x11xf32_1_1;
	end
	if (1'b1 == current_fsm_state06) begin
	    fadd_0_0_0_0_1_x <= fadd_0_0_0_0_1_r;
	    fadd_0_0_0_0_1_y <= fmul_0_0_0_0_1_r;
	end

	if (1'b1 == current_fsm_state07) begin
	    fmul_0_0_0_0_1_x <= p__arg0_0_2;
	    fmul_0_0_0_0_1_y <= p___constant_11x11xf32_1_2;
	end
	if (1'b1 == current_fsm_state09) begin
	    fadd_0_0_0_0_1_x <= fadd_0_0_0_0_1_r;
	    fadd_0_0_0_0_1_y <= fmul_0_0_0_0_1_r;
	end

	if (1'b1 == current_fsm_state10) begin
	    fmul_0_0_0_0_1_x <= p__arg0_0_3;
	    fmul_0_0_0_0_1_y <= p___constant_11x11xf32_1_3;
	end
	if (1'b1 == current_fsm_state12) begin
	    fadd_0_0_0_0_1_x <= fadd_0_0_0_0_1_r;
	    fadd_0_0_0_0_1_y <= fmul_0_0_0_0_1_r;
	end

	if (1'b1 == current_fsm_state13) begin
	    fmul_0_0_0_0_1_x <= p__arg0_0_4;
	    fmul_0_0_0_0_1_y <= p___constant_11x11xf32_1_4;
	end
	if (1'b1 == current_fsm_state15) begin
	    fadd_0_0_0_0_1_x <= fadd_0_0_0_0_1_r;
	    fadd_0_0_0_0_1_y <= fmul_0_0_0_0_1_r;
	end

	if (1'b1 == current_fsm_state16) begin
	    fmul_0_0_0_0_1_x <= p__arg0_0_5;
	    fmul_0_0_0_0_1_y <= p___constant_11x11xf32_1_5;
	end
	if (1'b1 == current_fsm_state18) begin
	    fadd_0_0_0_0_1_x <= fadd_0_0_0_0_1_r;
	    fadd_0_0_0_0_1_y <= fmul_0_0_0_0_1_r;
	end

	if (1'b1 == current_fsm_state19) begin
	    fmul_0_0_0_0_1_x <= p__arg0_0_6;
	    fmul_0_0_0_0_1_y <= p___constant_11x11xf32_1_6;
	end
	if (1'b1 == current_fsm_state21) begin
	    fadd_0_0_0_0_1_x <= fadd_0_0_0_0_1_r;
	    fadd_0_0_0_0_1_y <= fmul_0_0_0_0_1_r;
	end

	if (1'b1 == current_fsm_state22) begin
	    fmul_0_0_0_0_1_x <= p__arg0_0_7;
	    fmul_0_0_0_0_1_y <= p___constant_11x11xf32_1_7;
	end
	if (1'b1 == current_fsm_state24) begin
	    fadd_0_0_0_0_1_x <= fadd_0_0_0_0_1_r;
	    fadd_0_0_0_0_1_y <= fmul_0_0_0_0_1_r;
	end

	if (1'b1 == current_fsm_state25) begin
	    fmul_0_0_0_0_1_x <= p__arg0_0_8;
	    fmul_0_0_0_0_1_y <= p___constant_11x11xf32_1_8;
	end
	if (1'b1 == current_fsm_state27) begin
	    fadd_0_0_0_0_1_x <= fadd_0_0_0_0_1_r;
	    fadd_0_0_0_0_1_y <= fmul_0_0_0_0_1_r;
	end

	if (1'b1 == current_fsm_state28) begin
	    fmul_0_0_0_0_1_x <= p__arg0_0_9;
	    fmul_0_0_0_0_1_y <= p___constant_11x11xf32_1_9;
	end
	if (1'b1 == current_fsm_state30) begin
	    fadd_0_0_0_0_1_x <= fadd_0_0_0_0_1_r;
	    fadd_0_0_0_0_1_y <= fmul_0_0_0_0_1_r;
	end

	if (1'b1 == current_fsm_state31) begin
	    fmul_0_0_0_0_1_x <= p__arg0_0_10;
	    fmul_0_0_0_0_1_y <= p___constant_11x11xf32_1_10;
	end
	if (1'b1 == current_fsm_state33) begin
	    fadd_0_0_0_0_1_x <= fadd_0_0_0_0_1_r;
	    fadd_0_0_0_0_1_y <= fmul_0_0_0_0_1_r;
	end

	// p_val_58 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_1_0, p__arg0_0_1, p___constant_11x11xf32_1_1, p__arg0_0_2, p___constant_11x11xf32_1_2, p__arg0_0_3, p___constant_11x11xf32_1_3, p__arg0_0_4, p___constant_11x11xf32_1_4, p__arg0_0_5, p___constant_11x11xf32_1_5, p__arg0_0_6, p___constant_11x11xf32_1_6, p__arg0_0_7, p___constant_11x11xf32_1_7, p__arg0_0_8, p___constant_11x11xf32_1_8, p__arg0_0_9, p___constant_11x11xf32_1_9, p__arg0_0_10, p___constant_11x11xf32_1_10) {  pe = "(0, 0, 0, 0, 1)", opr = "fmac", op_id = "3", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 end


	// p_val_59 = "copy" (p_val_58) {  pe = "(0, 0, 0, 0, 1)", opr = "copy", op_id = "4", start_time = "36"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state36) begin
	    p_val_59 <= fadd_0_0_0_0_1_r;
	end
	// p_val_59 = "copy" (p_val_58) {  pe = "(0, 0, 0, 0, 1)", opr = "copy", op_id = "4", start_time = "36"  } : (f32) -> f32 end


	// p_val_277 = "fadd" (p_val_59, p___constant_11xf32_1) {  pe = "(0, 0, 0, 0, 1)", opr = "fadd", op_id = "24", start_time = "37"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state37) begin
	    fadd_0_0_0_0_1_x <= p_val_59;
	    fadd_0_0_0_0_1_y <= p___constant_11xf32_1;
	end
	// p_val_277 = "fadd" (p_val_59, p___constant_11xf32_1) {  pe = "(0, 0, 0, 0, 1)", opr = "fadd", op_id = "24", start_time = "37"  } : (f32, f32) -> f32 end


	// p_val_288 = "copy" (p_val_277) {  pe = "(0, 0, 0, 0, 1)", opr = "copy", op_id = "35", start_time = "40"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state40) begin
	    p_val_288 <= fadd_0_0_0_0_1_r;
	end
	// p_val_288 = "copy" (p_val_277) {  pe = "(0, 0, 0, 0, 1)", opr = "copy", op_id = "35", start_time = "40"  } : (f32) -> f32 end

end

always @ (posedge clk) begin

	// p_val_82 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_2_0, p__arg0_0_1, p___constant_11x11xf32_2_1, p__arg0_0_2, p___constant_11x11xf32_2_2, p__arg0_0_3, p___constant_11x11xf32_2_3, p__arg0_0_4, p___constant_11x11xf32_2_4, p__arg0_0_5, p___constant_11x11xf32_2_5, p__arg0_0_6, p___constant_11x11xf32_2_6, p__arg0_0_7, p___constant_11x11xf32_2_7, p__arg0_0_8, p___constant_11x11xf32_2_8, p__arg0_0_9, p___constant_11x11xf32_2_9, p__arg0_0_10, p___constant_11x11xf32_2_10) {  pe = "(0, 0, 0, 0, 2)", opr = "fmac", op_id = "5", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 start
	if (1'b1 == current_fsm_state01) begin
	    fmul_0_0_0_0_2_x <= p__arg0_0_0;
	    fmul_0_0_0_0_2_y <= p___constant_11x11xf32_2_0;
	end
	if (1'b1 == current_fsm_state03) begin
	    fadd_0_0_0_0_2_x <= p_val_cst_0_point_0000000000000000000000000;
	    fadd_0_0_0_0_2_y <= fmul_0_0_0_0_2_r;
	end

	if (1'b1 == current_fsm_state04) begin
	    fmul_0_0_0_0_2_x <= p__arg0_0_1;
	    fmul_0_0_0_0_2_y <= p___constant_11x11xf32_2_1;
	end
	if (1'b1 == current_fsm_state06) begin
	    fadd_0_0_0_0_2_x <= fadd_0_0_0_0_2_r;
	    fadd_0_0_0_0_2_y <= fmul_0_0_0_0_2_r;
	end

	if (1'b1 == current_fsm_state07) begin
	    fmul_0_0_0_0_2_x <= p__arg0_0_2;
	    fmul_0_0_0_0_2_y <= p___constant_11x11xf32_2_2;
	end
	if (1'b1 == current_fsm_state09) begin
	    fadd_0_0_0_0_2_x <= fadd_0_0_0_0_2_r;
	    fadd_0_0_0_0_2_y <= fmul_0_0_0_0_2_r;
	end

	if (1'b1 == current_fsm_state10) begin
	    fmul_0_0_0_0_2_x <= p__arg0_0_3;
	    fmul_0_0_0_0_2_y <= p___constant_11x11xf32_2_3;
	end
	if (1'b1 == current_fsm_state12) begin
	    fadd_0_0_0_0_2_x <= fadd_0_0_0_0_2_r;
	    fadd_0_0_0_0_2_y <= fmul_0_0_0_0_2_r;
	end

	if (1'b1 == current_fsm_state13) begin
	    fmul_0_0_0_0_2_x <= p__arg0_0_4;
	    fmul_0_0_0_0_2_y <= p___constant_11x11xf32_2_4;
	end
	if (1'b1 == current_fsm_state15) begin
	    fadd_0_0_0_0_2_x <= fadd_0_0_0_0_2_r;
	    fadd_0_0_0_0_2_y <= fmul_0_0_0_0_2_r;
	end

	if (1'b1 == current_fsm_state16) begin
	    fmul_0_0_0_0_2_x <= p__arg0_0_5;
	    fmul_0_0_0_0_2_y <= p___constant_11x11xf32_2_5;
	end
	if (1'b1 == current_fsm_state18) begin
	    fadd_0_0_0_0_2_x <= fadd_0_0_0_0_2_r;
	    fadd_0_0_0_0_2_y <= fmul_0_0_0_0_2_r;
	end

	if (1'b1 == current_fsm_state19) begin
	    fmul_0_0_0_0_2_x <= p__arg0_0_6;
	    fmul_0_0_0_0_2_y <= p___constant_11x11xf32_2_6;
	end
	if (1'b1 == current_fsm_state21) begin
	    fadd_0_0_0_0_2_x <= fadd_0_0_0_0_2_r;
	    fadd_0_0_0_0_2_y <= fmul_0_0_0_0_2_r;
	end

	if (1'b1 == current_fsm_state22) begin
	    fmul_0_0_0_0_2_x <= p__arg0_0_7;
	    fmul_0_0_0_0_2_y <= p___constant_11x11xf32_2_7;
	end
	if (1'b1 == current_fsm_state24) begin
	    fadd_0_0_0_0_2_x <= fadd_0_0_0_0_2_r;
	    fadd_0_0_0_0_2_y <= fmul_0_0_0_0_2_r;
	end

	if (1'b1 == current_fsm_state25) begin
	    fmul_0_0_0_0_2_x <= p__arg0_0_8;
	    fmul_0_0_0_0_2_y <= p___constant_11x11xf32_2_8;
	end
	if (1'b1 == current_fsm_state27) begin
	    fadd_0_0_0_0_2_x <= fadd_0_0_0_0_2_r;
	    fadd_0_0_0_0_2_y <= fmul_0_0_0_0_2_r;
	end

	if (1'b1 == current_fsm_state28) begin
	    fmul_0_0_0_0_2_x <= p__arg0_0_9;
	    fmul_0_0_0_0_2_y <= p___constant_11x11xf32_2_9;
	end
	if (1'b1 == current_fsm_state30) begin
	    fadd_0_0_0_0_2_x <= fadd_0_0_0_0_2_r;
	    fadd_0_0_0_0_2_y <= fmul_0_0_0_0_2_r;
	end

	if (1'b1 == current_fsm_state31) begin
	    fmul_0_0_0_0_2_x <= p__arg0_0_10;
	    fmul_0_0_0_0_2_y <= p___constant_11x11xf32_2_10;
	end
	if (1'b1 == current_fsm_state33) begin
	    fadd_0_0_0_0_2_x <= fadd_0_0_0_0_2_r;
	    fadd_0_0_0_0_2_y <= fmul_0_0_0_0_2_r;
	end

	// p_val_82 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_2_0, p__arg0_0_1, p___constant_11x11xf32_2_1, p__arg0_0_2, p___constant_11x11xf32_2_2, p__arg0_0_3, p___constant_11x11xf32_2_3, p__arg0_0_4, p___constant_11x11xf32_2_4, p__arg0_0_5, p___constant_11x11xf32_2_5, p__arg0_0_6, p___constant_11x11xf32_2_6, p__arg0_0_7, p___constant_11x11xf32_2_7, p__arg0_0_8, p___constant_11x11xf32_2_8, p__arg0_0_9, p___constant_11x11xf32_2_9, p__arg0_0_10, p___constant_11x11xf32_2_10) {  pe = "(0, 0, 0, 0, 2)", opr = "fmac", op_id = "5", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 end


	// p_val_83 = "copy" (p_val_82) {  pe = "(0, 0, 0, 0, 2)", opr = "copy", op_id = "6", start_time = "36"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state36) begin
	    p_val_83 <= fadd_0_0_0_0_2_r;
	end
	// p_val_83 = "copy" (p_val_82) {  pe = "(0, 0, 0, 0, 2)", opr = "copy", op_id = "6", start_time = "36"  } : (f32) -> f32 end


	// p_val_278 = "fadd" (p_val_83, p___constant_11xf32_2) {  pe = "(0, 0, 0, 0, 2)", opr = "fadd", op_id = "25", start_time = "37"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state37) begin
	    fadd_0_0_0_0_2_x <= p_val_83;
	    fadd_0_0_0_0_2_y <= p___constant_11xf32_2;
	end
	// p_val_278 = "fadd" (p_val_83, p___constant_11xf32_2) {  pe = "(0, 0, 0, 0, 2)", opr = "fadd", op_id = "25", start_time = "37"  } : (f32, f32) -> f32 end


	// p_val_289 = "copy" (p_val_278) {  pe = "(0, 0, 0, 0, 2)", opr = "copy", op_id = "36", start_time = "40"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state40) begin
	    p_val_289 <= fadd_0_0_0_0_2_r;
	end
	// p_val_289 = "copy" (p_val_278) {  pe = "(0, 0, 0, 0, 2)", opr = "copy", op_id = "36", start_time = "40"  } : (f32) -> f32 end


	// p_val_300 = "fadd" (p_val_289, p_val_290) {  pe = "(0, 0, 0, 0, 2)", opr = "fadd", op_id = "46", start_time = "41"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state41) begin
	    fadd_0_0_0_0_2_x <= p_val_289;
	    fadd_0_0_0_0_2_y <= p_val_290;
	end
	// p_val_300 = "fadd" (p_val_289, p_val_290) {  pe = "(0, 0, 0, 0, 2)", opr = "fadd", op_id = "46", start_time = "41"  } : (f32, f32) -> f32 end

end

always @ (posedge clk) begin

	// p_val_106 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_3_0, p__arg0_0_1, p___constant_11x11xf32_3_1, p__arg0_0_2, p___constant_11x11xf32_3_2, p__arg0_0_3, p___constant_11x11xf32_3_3, p__arg0_0_4, p___constant_11x11xf32_3_4, p__arg0_0_5, p___constant_11x11xf32_3_5, p__arg0_0_6, p___constant_11x11xf32_3_6, p__arg0_0_7, p___constant_11x11xf32_3_7, p__arg0_0_8, p___constant_11x11xf32_3_8, p__arg0_0_9, p___constant_11x11xf32_3_9, p__arg0_0_10, p___constant_11x11xf32_3_10) {  pe = "(0, 0, 0, 0, 3)", opr = "fmac", op_id = "7", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 start
	if (1'b1 == current_fsm_state01) begin
	    fmul_0_0_0_0_3_x <= p__arg0_0_0;
	    fmul_0_0_0_0_3_y <= p___constant_11x11xf32_3_0;
	end
	if (1'b1 == current_fsm_state03) begin
	    fadd_0_0_0_0_3_x <= p_val_cst_0_point_0000000000000000000000000;
	    fadd_0_0_0_0_3_y <= fmul_0_0_0_0_3_r;
	end

	if (1'b1 == current_fsm_state04) begin
	    fmul_0_0_0_0_3_x <= p__arg0_0_1;
	    fmul_0_0_0_0_3_y <= p___constant_11x11xf32_3_1;
	end
	if (1'b1 == current_fsm_state06) begin
	    fadd_0_0_0_0_3_x <= fadd_0_0_0_0_3_r;
	    fadd_0_0_0_0_3_y <= fmul_0_0_0_0_3_r;
	end

	if (1'b1 == current_fsm_state07) begin
	    fmul_0_0_0_0_3_x <= p__arg0_0_2;
	    fmul_0_0_0_0_3_y <= p___constant_11x11xf32_3_2;
	end
	if (1'b1 == current_fsm_state09) begin
	    fadd_0_0_0_0_3_x <= fadd_0_0_0_0_3_r;
	    fadd_0_0_0_0_3_y <= fmul_0_0_0_0_3_r;
	end

	if (1'b1 == current_fsm_state10) begin
	    fmul_0_0_0_0_3_x <= p__arg0_0_3;
	    fmul_0_0_0_0_3_y <= p___constant_11x11xf32_3_3;
	end
	if (1'b1 == current_fsm_state12) begin
	    fadd_0_0_0_0_3_x <= fadd_0_0_0_0_3_r;
	    fadd_0_0_0_0_3_y <= fmul_0_0_0_0_3_r;
	end

	if (1'b1 == current_fsm_state13) begin
	    fmul_0_0_0_0_3_x <= p__arg0_0_4;
	    fmul_0_0_0_0_3_y <= p___constant_11x11xf32_3_4;
	end
	if (1'b1 == current_fsm_state15) begin
	    fadd_0_0_0_0_3_x <= fadd_0_0_0_0_3_r;
	    fadd_0_0_0_0_3_y <= fmul_0_0_0_0_3_r;
	end

	if (1'b1 == current_fsm_state16) begin
	    fmul_0_0_0_0_3_x <= p__arg0_0_5;
	    fmul_0_0_0_0_3_y <= p___constant_11x11xf32_3_5;
	end
	if (1'b1 == current_fsm_state18) begin
	    fadd_0_0_0_0_3_x <= fadd_0_0_0_0_3_r;
	    fadd_0_0_0_0_3_y <= fmul_0_0_0_0_3_r;
	end

	if (1'b1 == current_fsm_state19) begin
	    fmul_0_0_0_0_3_x <= p__arg0_0_6;
	    fmul_0_0_0_0_3_y <= p___constant_11x11xf32_3_6;
	end
	if (1'b1 == current_fsm_state21) begin
	    fadd_0_0_0_0_3_x <= fadd_0_0_0_0_3_r;
	    fadd_0_0_0_0_3_y <= fmul_0_0_0_0_3_r;
	end

	if (1'b1 == current_fsm_state22) begin
	    fmul_0_0_0_0_3_x <= p__arg0_0_7;
	    fmul_0_0_0_0_3_y <= p___constant_11x11xf32_3_7;
	end
	if (1'b1 == current_fsm_state24) begin
	    fadd_0_0_0_0_3_x <= fadd_0_0_0_0_3_r;
	    fadd_0_0_0_0_3_y <= fmul_0_0_0_0_3_r;
	end

	if (1'b1 == current_fsm_state25) begin
	    fmul_0_0_0_0_3_x <= p__arg0_0_8;
	    fmul_0_0_0_0_3_y <= p___constant_11x11xf32_3_8;
	end
	if (1'b1 == current_fsm_state27) begin
	    fadd_0_0_0_0_3_x <= fadd_0_0_0_0_3_r;
	    fadd_0_0_0_0_3_y <= fmul_0_0_0_0_3_r;
	end

	if (1'b1 == current_fsm_state28) begin
	    fmul_0_0_0_0_3_x <= p__arg0_0_9;
	    fmul_0_0_0_0_3_y <= p___constant_11x11xf32_3_9;
	end
	if (1'b1 == current_fsm_state30) begin
	    fadd_0_0_0_0_3_x <= fadd_0_0_0_0_3_r;
	    fadd_0_0_0_0_3_y <= fmul_0_0_0_0_3_r;
	end

	if (1'b1 == current_fsm_state31) begin
	    fmul_0_0_0_0_3_x <= p__arg0_0_10;
	    fmul_0_0_0_0_3_y <= p___constant_11x11xf32_3_10;
	end
	if (1'b1 == current_fsm_state33) begin
	    fadd_0_0_0_0_3_x <= fadd_0_0_0_0_3_r;
	    fadd_0_0_0_0_3_y <= fmul_0_0_0_0_3_r;
	end

	// p_val_106 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_3_0, p__arg0_0_1, p___constant_11x11xf32_3_1, p__arg0_0_2, p___constant_11x11xf32_3_2, p__arg0_0_3, p___constant_11x11xf32_3_3, p__arg0_0_4, p___constant_11x11xf32_3_4, p__arg0_0_5, p___constant_11x11xf32_3_5, p__arg0_0_6, p___constant_11x11xf32_3_6, p__arg0_0_7, p___constant_11x11xf32_3_7, p__arg0_0_8, p___constant_11x11xf32_3_8, p__arg0_0_9, p___constant_11x11xf32_3_9, p__arg0_0_10, p___constant_11x11xf32_3_10) {  pe = "(0, 0, 0, 0, 3)", opr = "fmac", op_id = "7", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 end


	// p_val_107 = "copy" (p_val_106) {  pe = "(0, 0, 0, 0, 3)", opr = "copy", op_id = "8", start_time = "36"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state36) begin
	    p_val_107 <= fadd_0_0_0_0_3_r;
	end
	// p_val_107 = "copy" (p_val_106) {  pe = "(0, 0, 0, 0, 3)", opr = "copy", op_id = "8", start_time = "36"  } : (f32) -> f32 end


	// p_val_279 = "fadd" (p_val_107, p___constant_11xf32_3) {  pe = "(0, 0, 0, 0, 3)", opr = "fadd", op_id = "26", start_time = "37"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state37) begin
	    fadd_0_0_0_0_3_x <= p_val_107;
	    fadd_0_0_0_0_3_y <= p___constant_11xf32_3;
	end
	// p_val_279 = "fadd" (p_val_107, p___constant_11xf32_3) {  pe = "(0, 0, 0, 0, 3)", opr = "fadd", op_id = "26", start_time = "37"  } : (f32, f32) -> f32 end


	// p_val_290 = "copy" (p_val_279) {  pe = "(0, 0, 0, 0, 3)", opr = "copy", op_id = "37", start_time = "40"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state40) begin
	    p_val_290 <= fadd_0_0_0_0_3_r;
	end
	// p_val_290 = "copy" (p_val_279) {  pe = "(0, 0, 0, 0, 3)", opr = "copy", op_id = "37", start_time = "40"  } : (f32) -> f32 end

end

always @ (posedge clk) begin

	// p_val_130 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_4_0, p__arg0_0_1, p___constant_11x11xf32_4_1, p__arg0_0_2, p___constant_11x11xf32_4_2, p__arg0_0_3, p___constant_11x11xf32_4_3, p__arg0_0_4, p___constant_11x11xf32_4_4, p__arg0_0_5, p___constant_11x11xf32_4_5, p__arg0_0_6, p___constant_11x11xf32_4_6, p__arg0_0_7, p___constant_11x11xf32_4_7, p__arg0_0_8, p___constant_11x11xf32_4_8, p__arg0_0_9, p___constant_11x11xf32_4_9, p__arg0_0_10, p___constant_11x11xf32_4_10) {  pe = "(0, 0, 0, 0, 4)", opr = "fmac", op_id = "9", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 start
	if (1'b1 == current_fsm_state01) begin
	    fmul_0_0_0_0_4_x <= p__arg0_0_0;
	    fmul_0_0_0_0_4_y <= p___constant_11x11xf32_4_0;
	end
	if (1'b1 == current_fsm_state03) begin
	    fadd_0_0_0_0_4_x <= p_val_cst_0_point_0000000000000000000000000;
	    fadd_0_0_0_0_4_y <= fmul_0_0_0_0_4_r;
	end

	if (1'b1 == current_fsm_state04) begin
	    fmul_0_0_0_0_4_x <= p__arg0_0_1;
	    fmul_0_0_0_0_4_y <= p___constant_11x11xf32_4_1;
	end
	if (1'b1 == current_fsm_state06) begin
	    fadd_0_0_0_0_4_x <= fadd_0_0_0_0_4_r;
	    fadd_0_0_0_0_4_y <= fmul_0_0_0_0_4_r;
	end

	if (1'b1 == current_fsm_state07) begin
	    fmul_0_0_0_0_4_x <= p__arg0_0_2;
	    fmul_0_0_0_0_4_y <= p___constant_11x11xf32_4_2;
	end
	if (1'b1 == current_fsm_state09) begin
	    fadd_0_0_0_0_4_x <= fadd_0_0_0_0_4_r;
	    fadd_0_0_0_0_4_y <= fmul_0_0_0_0_4_r;
	end

	if (1'b1 == current_fsm_state10) begin
	    fmul_0_0_0_0_4_x <= p__arg0_0_3;
	    fmul_0_0_0_0_4_y <= p___constant_11x11xf32_4_3;
	end
	if (1'b1 == current_fsm_state12) begin
	    fadd_0_0_0_0_4_x <= fadd_0_0_0_0_4_r;
	    fadd_0_0_0_0_4_y <= fmul_0_0_0_0_4_r;
	end

	if (1'b1 == current_fsm_state13) begin
	    fmul_0_0_0_0_4_x <= p__arg0_0_4;
	    fmul_0_0_0_0_4_y <= p___constant_11x11xf32_4_4;
	end
	if (1'b1 == current_fsm_state15) begin
	    fadd_0_0_0_0_4_x <= fadd_0_0_0_0_4_r;
	    fadd_0_0_0_0_4_y <= fmul_0_0_0_0_4_r;
	end

	if (1'b1 == current_fsm_state16) begin
	    fmul_0_0_0_0_4_x <= p__arg0_0_5;
	    fmul_0_0_0_0_4_y <= p___constant_11x11xf32_4_5;
	end
	if (1'b1 == current_fsm_state18) begin
	    fadd_0_0_0_0_4_x <= fadd_0_0_0_0_4_r;
	    fadd_0_0_0_0_4_y <= fmul_0_0_0_0_4_r;
	end

	if (1'b1 == current_fsm_state19) begin
	    fmul_0_0_0_0_4_x <= p__arg0_0_6;
	    fmul_0_0_0_0_4_y <= p___constant_11x11xf32_4_6;
	end
	if (1'b1 == current_fsm_state21) begin
	    fadd_0_0_0_0_4_x <= fadd_0_0_0_0_4_r;
	    fadd_0_0_0_0_4_y <= fmul_0_0_0_0_4_r;
	end

	if (1'b1 == current_fsm_state22) begin
	    fmul_0_0_0_0_4_x <= p__arg0_0_7;
	    fmul_0_0_0_0_4_y <= p___constant_11x11xf32_4_7;
	end
	if (1'b1 == current_fsm_state24) begin
	    fadd_0_0_0_0_4_x <= fadd_0_0_0_0_4_r;
	    fadd_0_0_0_0_4_y <= fmul_0_0_0_0_4_r;
	end

	if (1'b1 == current_fsm_state25) begin
	    fmul_0_0_0_0_4_x <= p__arg0_0_8;
	    fmul_0_0_0_0_4_y <= p___constant_11x11xf32_4_8;
	end
	if (1'b1 == current_fsm_state27) begin
	    fadd_0_0_0_0_4_x <= fadd_0_0_0_0_4_r;
	    fadd_0_0_0_0_4_y <= fmul_0_0_0_0_4_r;
	end

	if (1'b1 == current_fsm_state28) begin
	    fmul_0_0_0_0_4_x <= p__arg0_0_9;
	    fmul_0_0_0_0_4_y <= p___constant_11x11xf32_4_9;
	end
	if (1'b1 == current_fsm_state30) begin
	    fadd_0_0_0_0_4_x <= fadd_0_0_0_0_4_r;
	    fadd_0_0_0_0_4_y <= fmul_0_0_0_0_4_r;
	end

	if (1'b1 == current_fsm_state31) begin
	    fmul_0_0_0_0_4_x <= p__arg0_0_10;
	    fmul_0_0_0_0_4_y <= p___constant_11x11xf32_4_10;
	end
	if (1'b1 == current_fsm_state33) begin
	    fadd_0_0_0_0_4_x <= fadd_0_0_0_0_4_r;
	    fadd_0_0_0_0_4_y <= fmul_0_0_0_0_4_r;
	end

	// p_val_130 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_4_0, p__arg0_0_1, p___constant_11x11xf32_4_1, p__arg0_0_2, p___constant_11x11xf32_4_2, p__arg0_0_3, p___constant_11x11xf32_4_3, p__arg0_0_4, p___constant_11x11xf32_4_4, p__arg0_0_5, p___constant_11x11xf32_4_5, p__arg0_0_6, p___constant_11x11xf32_4_6, p__arg0_0_7, p___constant_11x11xf32_4_7, p__arg0_0_8, p___constant_11x11xf32_4_8, p__arg0_0_9, p___constant_11x11xf32_4_9, p__arg0_0_10, p___constant_11x11xf32_4_10) {  pe = "(0, 0, 0, 0, 4)", opr = "fmac", op_id = "9", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 end


	// p_val_131 = "copy" (p_val_130) {  pe = "(0, 0, 0, 0, 4)", opr = "copy", op_id = "10", start_time = "36"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state36) begin
	    p_val_131 <= fadd_0_0_0_0_4_r;
	end
	// p_val_131 = "copy" (p_val_130) {  pe = "(0, 0, 0, 0, 4)", opr = "copy", op_id = "10", start_time = "36"  } : (f32) -> f32 end


	// p_val_280 = "fadd" (p_val_131, p___constant_11xf32_4) {  pe = "(0, 0, 0, 0, 4)", opr = "fadd", op_id = "27", start_time = "37"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state37) begin
	    fadd_0_0_0_0_4_x <= p_val_131;
	    fadd_0_0_0_0_4_y <= p___constant_11xf32_4;
	end
	// p_val_280 = "fadd" (p_val_131, p___constant_11xf32_4) {  pe = "(0, 0, 0, 0, 4)", opr = "fadd", op_id = "27", start_time = "37"  } : (f32, f32) -> f32 end


	// p_val_291 = "copy" (p_val_280) {  pe = "(0, 0, 0, 0, 4)", opr = "copy", op_id = "38", start_time = "40"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state40) begin
	    p_val_291 <= fadd_0_0_0_0_4_r;
	end
	// p_val_291 = "copy" (p_val_280) {  pe = "(0, 0, 0, 0, 4)", opr = "copy", op_id = "38", start_time = "40"  } : (f32) -> f32 end


	// p_val_301 = "fadd" (p_val_291, p_val_292) {  pe = "(0, 0, 0, 0, 4)", opr = "fadd", op_id = "47", start_time = "41"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state41) begin
	    fadd_0_0_0_0_4_x <= p_val_291;
	    fadd_0_0_0_0_4_y <= p_val_292;
	end
	// p_val_301 = "fadd" (p_val_291, p_val_292) {  pe = "(0, 0, 0, 0, 4)", opr = "fadd", op_id = "47", start_time = "41"  } : (f32, f32) -> f32 end


	// p_val_304 = "fadd" (p_val_301, p_val_302) {  pe = "(0, 0, 0, 0, 4)", opr = "fadd", op_id = "50", start_time = "44"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state44) begin
	    fadd_0_0_0_0_4_x <= fadd_0_0_0_0_4_r;
	    fadd_0_0_0_0_4_y <= fadd_0_0_0_0_6_r;
	end
	// p_val_304 = "fadd" (p_val_301, p_val_302) {  pe = "(0, 0, 0, 0, 4)", opr = "fadd", op_id = "50", start_time = "44"  } : (f32, f32) -> f32 end

end

always @ (posedge clk) begin

	// p_val_154 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_5_0, p__arg0_0_1, p___constant_11x11xf32_5_1, p__arg0_0_2, p___constant_11x11xf32_5_2, p__arg0_0_3, p___constant_11x11xf32_5_3, p__arg0_0_4, p___constant_11x11xf32_5_4, p__arg0_0_5, p___constant_11x11xf32_5_5, p__arg0_0_6, p___constant_11x11xf32_5_6, p__arg0_0_7, p___constant_11x11xf32_5_7, p__arg0_0_8, p___constant_11x11xf32_5_8, p__arg0_0_9, p___constant_11x11xf32_5_9, p__arg0_0_10, p___constant_11x11xf32_5_10) {  pe = "(0, 0, 0, 0, 5)", opr = "fmac", op_id = "11", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 start
	if (1'b1 == current_fsm_state01) begin
	    fmul_0_0_0_0_5_x <= p__arg0_0_0;
	    fmul_0_0_0_0_5_y <= p___constant_11x11xf32_5_0;
	end
	if (1'b1 == current_fsm_state03) begin
	    fadd_0_0_0_0_5_x <= p_val_cst_0_point_0000000000000000000000000;
	    fadd_0_0_0_0_5_y <= fmul_0_0_0_0_5_r;
	end

	if (1'b1 == current_fsm_state04) begin
	    fmul_0_0_0_0_5_x <= p__arg0_0_1;
	    fmul_0_0_0_0_5_y <= p___constant_11x11xf32_5_1;
	end
	if (1'b1 == current_fsm_state06) begin
	    fadd_0_0_0_0_5_x <= fadd_0_0_0_0_5_r;
	    fadd_0_0_0_0_5_y <= fmul_0_0_0_0_5_r;
	end

	if (1'b1 == current_fsm_state07) begin
	    fmul_0_0_0_0_5_x <= p__arg0_0_2;
	    fmul_0_0_0_0_5_y <= p___constant_11x11xf32_5_2;
	end
	if (1'b1 == current_fsm_state09) begin
	    fadd_0_0_0_0_5_x <= fadd_0_0_0_0_5_r;
	    fadd_0_0_0_0_5_y <= fmul_0_0_0_0_5_r;
	end

	if (1'b1 == current_fsm_state10) begin
	    fmul_0_0_0_0_5_x <= p__arg0_0_3;
	    fmul_0_0_0_0_5_y <= p___constant_11x11xf32_5_3;
	end
	if (1'b1 == current_fsm_state12) begin
	    fadd_0_0_0_0_5_x <= fadd_0_0_0_0_5_r;
	    fadd_0_0_0_0_5_y <= fmul_0_0_0_0_5_r;
	end

	if (1'b1 == current_fsm_state13) begin
	    fmul_0_0_0_0_5_x <= p__arg0_0_4;
	    fmul_0_0_0_0_5_y <= p___constant_11x11xf32_5_4;
	end
	if (1'b1 == current_fsm_state15) begin
	    fadd_0_0_0_0_5_x <= fadd_0_0_0_0_5_r;
	    fadd_0_0_0_0_5_y <= fmul_0_0_0_0_5_r;
	end

	if (1'b1 == current_fsm_state16) begin
	    fmul_0_0_0_0_5_x <= p__arg0_0_5;
	    fmul_0_0_0_0_5_y <= p___constant_11x11xf32_5_5;
	end
	if (1'b1 == current_fsm_state18) begin
	    fadd_0_0_0_0_5_x <= fadd_0_0_0_0_5_r;
	    fadd_0_0_0_0_5_y <= fmul_0_0_0_0_5_r;
	end

	if (1'b1 == current_fsm_state19) begin
	    fmul_0_0_0_0_5_x <= p__arg0_0_6;
	    fmul_0_0_0_0_5_y <= p___constant_11x11xf32_5_6;
	end
	if (1'b1 == current_fsm_state21) begin
	    fadd_0_0_0_0_5_x <= fadd_0_0_0_0_5_r;
	    fadd_0_0_0_0_5_y <= fmul_0_0_0_0_5_r;
	end

	if (1'b1 == current_fsm_state22) begin
	    fmul_0_0_0_0_5_x <= p__arg0_0_7;
	    fmul_0_0_0_0_5_y <= p___constant_11x11xf32_5_7;
	end
	if (1'b1 == current_fsm_state24) begin
	    fadd_0_0_0_0_5_x <= fadd_0_0_0_0_5_r;
	    fadd_0_0_0_0_5_y <= fmul_0_0_0_0_5_r;
	end

	if (1'b1 == current_fsm_state25) begin
	    fmul_0_0_0_0_5_x <= p__arg0_0_8;
	    fmul_0_0_0_0_5_y <= p___constant_11x11xf32_5_8;
	end
	if (1'b1 == current_fsm_state27) begin
	    fadd_0_0_0_0_5_x <= fadd_0_0_0_0_5_r;
	    fadd_0_0_0_0_5_y <= fmul_0_0_0_0_5_r;
	end

	if (1'b1 == current_fsm_state28) begin
	    fmul_0_0_0_0_5_x <= p__arg0_0_9;
	    fmul_0_0_0_0_5_y <= p___constant_11x11xf32_5_9;
	end
	if (1'b1 == current_fsm_state30) begin
	    fadd_0_0_0_0_5_x <= fadd_0_0_0_0_5_r;
	    fadd_0_0_0_0_5_y <= fmul_0_0_0_0_5_r;
	end

	if (1'b1 == current_fsm_state31) begin
	    fmul_0_0_0_0_5_x <= p__arg0_0_10;
	    fmul_0_0_0_0_5_y <= p___constant_11x11xf32_5_10;
	end
	if (1'b1 == current_fsm_state33) begin
	    fadd_0_0_0_0_5_x <= fadd_0_0_0_0_5_r;
	    fadd_0_0_0_0_5_y <= fmul_0_0_0_0_5_r;
	end

	// p_val_154 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_5_0, p__arg0_0_1, p___constant_11x11xf32_5_1, p__arg0_0_2, p___constant_11x11xf32_5_2, p__arg0_0_3, p___constant_11x11xf32_5_3, p__arg0_0_4, p___constant_11x11xf32_5_4, p__arg0_0_5, p___constant_11x11xf32_5_5, p__arg0_0_6, p___constant_11x11xf32_5_6, p__arg0_0_7, p___constant_11x11xf32_5_7, p__arg0_0_8, p___constant_11x11xf32_5_8, p__arg0_0_9, p___constant_11x11xf32_5_9, p__arg0_0_10, p___constant_11x11xf32_5_10) {  pe = "(0, 0, 0, 0, 5)", opr = "fmac", op_id = "11", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 end


	// p_val_155 = "copy" (p_val_154) {  pe = "(0, 0, 0, 0, 5)", opr = "copy", op_id = "12", start_time = "36"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state36) begin
	    p_val_155 <= fadd_0_0_0_0_5_r;
	end
	// p_val_155 = "copy" (p_val_154) {  pe = "(0, 0, 0, 0, 5)", opr = "copy", op_id = "12", start_time = "36"  } : (f32) -> f32 end


	// p_val_281 = "fadd" (p_val_155, p___constant_11xf32_5) {  pe = "(0, 0, 0, 0, 5)", opr = "fadd", op_id = "28", start_time = "37"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state37) begin
	    fadd_0_0_0_0_5_x <= p_val_155;
	    fadd_0_0_0_0_5_y <= p___constant_11xf32_5;
	end
	// p_val_281 = "fadd" (p_val_155, p___constant_11xf32_5) {  pe = "(0, 0, 0, 0, 5)", opr = "fadd", op_id = "28", start_time = "37"  } : (f32, f32) -> f32 end


	// p_val_292 = "copy" (p_val_281) {  pe = "(0, 0, 0, 0, 5)", opr = "copy", op_id = "39", start_time = "40"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state40) begin
	    p_val_292 <= fadd_0_0_0_0_5_r;
	end
	// p_val_292 = "copy" (p_val_281) {  pe = "(0, 0, 0, 0, 5)", opr = "copy", op_id = "39", start_time = "40"  } : (f32) -> f32 end

end

always @ (posedge clk) begin

	// p_val_178 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_6_0, p__arg0_0_1, p___constant_11x11xf32_6_1, p__arg0_0_2, p___constant_11x11xf32_6_2, p__arg0_0_3, p___constant_11x11xf32_6_3, p__arg0_0_4, p___constant_11x11xf32_6_4, p__arg0_0_5, p___constant_11x11xf32_6_5, p__arg0_0_6, p___constant_11x11xf32_6_6, p__arg0_0_7, p___constant_11x11xf32_6_7, p__arg0_0_8, p___constant_11x11xf32_6_8, p__arg0_0_9, p___constant_11x11xf32_6_9, p__arg0_0_10, p___constant_11x11xf32_6_10) {  pe = "(0, 0, 0, 0, 6)", opr = "fmac", op_id = "13", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 start
	if (1'b1 == current_fsm_state01) begin
	    fmul_0_0_0_0_6_x <= p__arg0_0_0;
	    fmul_0_0_0_0_6_y <= p___constant_11x11xf32_6_0;
	end
	if (1'b1 == current_fsm_state03) begin
	    fadd_0_0_0_0_6_x <= p_val_cst_0_point_0000000000000000000000000;
	    fadd_0_0_0_0_6_y <= fmul_0_0_0_0_6_r;
	end

	if (1'b1 == current_fsm_state04) begin
	    fmul_0_0_0_0_6_x <= p__arg0_0_1;
	    fmul_0_0_0_0_6_y <= p___constant_11x11xf32_6_1;
	end
	if (1'b1 == current_fsm_state06) begin
	    fadd_0_0_0_0_6_x <= fadd_0_0_0_0_6_r;
	    fadd_0_0_0_0_6_y <= fmul_0_0_0_0_6_r;
	end

	if (1'b1 == current_fsm_state07) begin
	    fmul_0_0_0_0_6_x <= p__arg0_0_2;
	    fmul_0_0_0_0_6_y <= p___constant_11x11xf32_6_2;
	end
	if (1'b1 == current_fsm_state09) begin
	    fadd_0_0_0_0_6_x <= fadd_0_0_0_0_6_r;
	    fadd_0_0_0_0_6_y <= fmul_0_0_0_0_6_r;
	end

	if (1'b1 == current_fsm_state10) begin
	    fmul_0_0_0_0_6_x <= p__arg0_0_3;
	    fmul_0_0_0_0_6_y <= p___constant_11x11xf32_6_3;
	end
	if (1'b1 == current_fsm_state12) begin
	    fadd_0_0_0_0_6_x <= fadd_0_0_0_0_6_r;
	    fadd_0_0_0_0_6_y <= fmul_0_0_0_0_6_r;
	end

	if (1'b1 == current_fsm_state13) begin
	    fmul_0_0_0_0_6_x <= p__arg0_0_4;
	    fmul_0_0_0_0_6_y <= p___constant_11x11xf32_6_4;
	end
	if (1'b1 == current_fsm_state15) begin
	    fadd_0_0_0_0_6_x <= fadd_0_0_0_0_6_r;
	    fadd_0_0_0_0_6_y <= fmul_0_0_0_0_6_r;
	end

	if (1'b1 == current_fsm_state16) begin
	    fmul_0_0_0_0_6_x <= p__arg0_0_5;
	    fmul_0_0_0_0_6_y <= p___constant_11x11xf32_6_5;
	end
	if (1'b1 == current_fsm_state18) begin
	    fadd_0_0_0_0_6_x <= fadd_0_0_0_0_6_r;
	    fadd_0_0_0_0_6_y <= fmul_0_0_0_0_6_r;
	end

	if (1'b1 == current_fsm_state19) begin
	    fmul_0_0_0_0_6_x <= p__arg0_0_6;
	    fmul_0_0_0_0_6_y <= p___constant_11x11xf32_6_6;
	end
	if (1'b1 == current_fsm_state21) begin
	    fadd_0_0_0_0_6_x <= fadd_0_0_0_0_6_r;
	    fadd_0_0_0_0_6_y <= fmul_0_0_0_0_6_r;
	end

	if (1'b1 == current_fsm_state22) begin
	    fmul_0_0_0_0_6_x <= p__arg0_0_7;
	    fmul_0_0_0_0_6_y <= p___constant_11x11xf32_6_7;
	end
	if (1'b1 == current_fsm_state24) begin
	    fadd_0_0_0_0_6_x <= fadd_0_0_0_0_6_r;
	    fadd_0_0_0_0_6_y <= fmul_0_0_0_0_6_r;
	end

	if (1'b1 == current_fsm_state25) begin
	    fmul_0_0_0_0_6_x <= p__arg0_0_8;
	    fmul_0_0_0_0_6_y <= p___constant_11x11xf32_6_8;
	end
	if (1'b1 == current_fsm_state27) begin
	    fadd_0_0_0_0_6_x <= fadd_0_0_0_0_6_r;
	    fadd_0_0_0_0_6_y <= fmul_0_0_0_0_6_r;
	end

	if (1'b1 == current_fsm_state28) begin
	    fmul_0_0_0_0_6_x <= p__arg0_0_9;
	    fmul_0_0_0_0_6_y <= p___constant_11x11xf32_6_9;
	end
	if (1'b1 == current_fsm_state30) begin
	    fadd_0_0_0_0_6_x <= fadd_0_0_0_0_6_r;
	    fadd_0_0_0_0_6_y <= fmul_0_0_0_0_6_r;
	end

	if (1'b1 == current_fsm_state31) begin
	    fmul_0_0_0_0_6_x <= p__arg0_0_10;
	    fmul_0_0_0_0_6_y <= p___constant_11x11xf32_6_10;
	end
	if (1'b1 == current_fsm_state33) begin
	    fadd_0_0_0_0_6_x <= fadd_0_0_0_0_6_r;
	    fadd_0_0_0_0_6_y <= fmul_0_0_0_0_6_r;
	end

	// p_val_178 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_6_0, p__arg0_0_1, p___constant_11x11xf32_6_1, p__arg0_0_2, p___constant_11x11xf32_6_2, p__arg0_0_3, p___constant_11x11xf32_6_3, p__arg0_0_4, p___constant_11x11xf32_6_4, p__arg0_0_5, p___constant_11x11xf32_6_5, p__arg0_0_6, p___constant_11x11xf32_6_6, p__arg0_0_7, p___constant_11x11xf32_6_7, p__arg0_0_8, p___constant_11x11xf32_6_8, p__arg0_0_9, p___constant_11x11xf32_6_9, p__arg0_0_10, p___constant_11x11xf32_6_10) {  pe = "(0, 0, 0, 0, 6)", opr = "fmac", op_id = "13", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 end


	// p_val_179 = "copy" (p_val_178) {  pe = "(0, 0, 0, 0, 6)", opr = "copy", op_id = "14", start_time = "36"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state36) begin
	    p_val_179 <= fadd_0_0_0_0_6_r;
	end
	// p_val_179 = "copy" (p_val_178) {  pe = "(0, 0, 0, 0, 6)", opr = "copy", op_id = "14", start_time = "36"  } : (f32) -> f32 end


	// p_val_282 = "fadd" (p_val_179, p___constant_11xf32_6) {  pe = "(0, 0, 0, 0, 6)", opr = "fadd", op_id = "29", start_time = "37"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state37) begin
	    fadd_0_0_0_0_6_x <= p_val_179;
	    fadd_0_0_0_0_6_y <= p___constant_11xf32_6;
	end
	// p_val_282 = "fadd" (p_val_179, p___constant_11xf32_6) {  pe = "(0, 0, 0, 0, 6)", opr = "fadd", op_id = "29", start_time = "37"  } : (f32, f32) -> f32 end


	// p_val_293 = "copy" (p_val_282) {  pe = "(0, 0, 0, 0, 6)", opr = "copy", op_id = "40", start_time = "40"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state40) begin
	    p_val_293 <= fadd_0_0_0_0_6_r;
	end
	// p_val_293 = "copy" (p_val_282) {  pe = "(0, 0, 0, 0, 6)", opr = "copy", op_id = "40", start_time = "40"  } : (f32) -> f32 end


	// p_val_302 = "fadd" (p_val_293, p_val_294) {  pe = "(0, 0, 0, 0, 6)", opr = "fadd", op_id = "48", start_time = "41"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state41) begin
	    fadd_0_0_0_0_6_x <= p_val_293;
	    fadd_0_0_0_0_6_y <= p_val_294;
	end
	// p_val_302 = "fadd" (p_val_293, p_val_294) {  pe = "(0, 0, 0, 0, 6)", opr = "fadd", op_id = "48", start_time = "41"  } : (f32, f32) -> f32 end

end

always @ (posedge clk) begin

	// p_val_202 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_7_0, p__arg0_0_1, p___constant_11x11xf32_7_1, p__arg0_0_2, p___constant_11x11xf32_7_2, p__arg0_0_3, p___constant_11x11xf32_7_3, p__arg0_0_4, p___constant_11x11xf32_7_4, p__arg0_0_5, p___constant_11x11xf32_7_5, p__arg0_0_6, p___constant_11x11xf32_7_6, p__arg0_0_7, p___constant_11x11xf32_7_7, p__arg0_0_8, p___constant_11x11xf32_7_8, p__arg0_0_9, p___constant_11x11xf32_7_9, p__arg0_0_10, p___constant_11x11xf32_7_10) {  pe = "(0, 0, 0, 0, 7)", opr = "fmac", op_id = "15", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 start
	if (1'b1 == current_fsm_state01) begin
	    fmul_0_0_0_0_7_x <= p__arg0_0_0;
	    fmul_0_0_0_0_7_y <= p___constant_11x11xf32_7_0;
	end
	if (1'b1 == current_fsm_state03) begin
	    fadd_0_0_0_0_7_x <= p_val_cst_0_point_0000000000000000000000000;
	    fadd_0_0_0_0_7_y <= fmul_0_0_0_0_7_r;
	end

	if (1'b1 == current_fsm_state04) begin
	    fmul_0_0_0_0_7_x <= p__arg0_0_1;
	    fmul_0_0_0_0_7_y <= p___constant_11x11xf32_7_1;
	end
	if (1'b1 == current_fsm_state06) begin
	    fadd_0_0_0_0_7_x <= fadd_0_0_0_0_7_r;
	    fadd_0_0_0_0_7_y <= fmul_0_0_0_0_7_r;
	end

	if (1'b1 == current_fsm_state07) begin
	    fmul_0_0_0_0_7_x <= p__arg0_0_2;
	    fmul_0_0_0_0_7_y <= p___constant_11x11xf32_7_2;
	end
	if (1'b1 == current_fsm_state09) begin
	    fadd_0_0_0_0_7_x <= fadd_0_0_0_0_7_r;
	    fadd_0_0_0_0_7_y <= fmul_0_0_0_0_7_r;
	end

	if (1'b1 == current_fsm_state10) begin
	    fmul_0_0_0_0_7_x <= p__arg0_0_3;
	    fmul_0_0_0_0_7_y <= p___constant_11x11xf32_7_3;
	end
	if (1'b1 == current_fsm_state12) begin
	    fadd_0_0_0_0_7_x <= fadd_0_0_0_0_7_r;
	    fadd_0_0_0_0_7_y <= fmul_0_0_0_0_7_r;
	end

	if (1'b1 == current_fsm_state13) begin
	    fmul_0_0_0_0_7_x <= p__arg0_0_4;
	    fmul_0_0_0_0_7_y <= p___constant_11x11xf32_7_4;
	end
	if (1'b1 == current_fsm_state15) begin
	    fadd_0_0_0_0_7_x <= fadd_0_0_0_0_7_r;
	    fadd_0_0_0_0_7_y <= fmul_0_0_0_0_7_r;
	end

	if (1'b1 == current_fsm_state16) begin
	    fmul_0_0_0_0_7_x <= p__arg0_0_5;
	    fmul_0_0_0_0_7_y <= p___constant_11x11xf32_7_5;
	end
	if (1'b1 == current_fsm_state18) begin
	    fadd_0_0_0_0_7_x <= fadd_0_0_0_0_7_r;
	    fadd_0_0_0_0_7_y <= fmul_0_0_0_0_7_r;
	end

	if (1'b1 == current_fsm_state19) begin
	    fmul_0_0_0_0_7_x <= p__arg0_0_6;
	    fmul_0_0_0_0_7_y <= p___constant_11x11xf32_7_6;
	end
	if (1'b1 == current_fsm_state21) begin
	    fadd_0_0_0_0_7_x <= fadd_0_0_0_0_7_r;
	    fadd_0_0_0_0_7_y <= fmul_0_0_0_0_7_r;
	end

	if (1'b1 == current_fsm_state22) begin
	    fmul_0_0_0_0_7_x <= p__arg0_0_7;
	    fmul_0_0_0_0_7_y <= p___constant_11x11xf32_7_7;
	end
	if (1'b1 == current_fsm_state24) begin
	    fadd_0_0_0_0_7_x <= fadd_0_0_0_0_7_r;
	    fadd_0_0_0_0_7_y <= fmul_0_0_0_0_7_r;
	end

	if (1'b1 == current_fsm_state25) begin
	    fmul_0_0_0_0_7_x <= p__arg0_0_8;
	    fmul_0_0_0_0_7_y <= p___constant_11x11xf32_7_8;
	end
	if (1'b1 == current_fsm_state27) begin
	    fadd_0_0_0_0_7_x <= fadd_0_0_0_0_7_r;
	    fadd_0_0_0_0_7_y <= fmul_0_0_0_0_7_r;
	end

	if (1'b1 == current_fsm_state28) begin
	    fmul_0_0_0_0_7_x <= p__arg0_0_9;
	    fmul_0_0_0_0_7_y <= p___constant_11x11xf32_7_9;
	end
	if (1'b1 == current_fsm_state30) begin
	    fadd_0_0_0_0_7_x <= fadd_0_0_0_0_7_r;
	    fadd_0_0_0_0_7_y <= fmul_0_0_0_0_7_r;
	end

	if (1'b1 == current_fsm_state31) begin
	    fmul_0_0_0_0_7_x <= p__arg0_0_10;
	    fmul_0_0_0_0_7_y <= p___constant_11x11xf32_7_10;
	end
	if (1'b1 == current_fsm_state33) begin
	    fadd_0_0_0_0_7_x <= fadd_0_0_0_0_7_r;
	    fadd_0_0_0_0_7_y <= fmul_0_0_0_0_7_r;
	end

	// p_val_202 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_7_0, p__arg0_0_1, p___constant_11x11xf32_7_1, p__arg0_0_2, p___constant_11x11xf32_7_2, p__arg0_0_3, p___constant_11x11xf32_7_3, p__arg0_0_4, p___constant_11x11xf32_7_4, p__arg0_0_5, p___constant_11x11xf32_7_5, p__arg0_0_6, p___constant_11x11xf32_7_6, p__arg0_0_7, p___constant_11x11xf32_7_7, p__arg0_0_8, p___constant_11x11xf32_7_8, p__arg0_0_9, p___constant_11x11xf32_7_9, p__arg0_0_10, p___constant_11x11xf32_7_10) {  pe = "(0, 0, 0, 0, 7)", opr = "fmac", op_id = "15", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 end


	// p_val_203 = "copy" (p_val_202) {  pe = "(0, 0, 0, 0, 7)", opr = "copy", op_id = "16", start_time = "36"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state36) begin
	    p_val_203 <= fadd_0_0_0_0_7_r;
	end
	// p_val_203 = "copy" (p_val_202) {  pe = "(0, 0, 0, 0, 7)", opr = "copy", op_id = "16", start_time = "36"  } : (f32) -> f32 end


	// p_val_283 = "fadd" (p_val_203, p___constant_11xf32_7) {  pe = "(0, 0, 0, 0, 7)", opr = "fadd", op_id = "30", start_time = "37"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state37) begin
	    fadd_0_0_0_0_7_x <= p_val_203;
	    fadd_0_0_0_0_7_y <= p___constant_11xf32_7;
	end
	// p_val_283 = "fadd" (p_val_203, p___constant_11xf32_7) {  pe = "(0, 0, 0, 0, 7)", opr = "fadd", op_id = "30", start_time = "37"  } : (f32, f32) -> f32 end


	// p_val_294 = "copy" (p_val_283) {  pe = "(0, 0, 0, 0, 7)", opr = "copy", op_id = "41", start_time = "40"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state40) begin
	    p_val_294 <= fadd_0_0_0_0_7_r;
	end
	// p_val_294 = "copy" (p_val_283) {  pe = "(0, 0, 0, 0, 7)", opr = "copy", op_id = "41", start_time = "40"  } : (f32) -> f32 end

end

always @ (posedge clk) begin

	// p_val_226 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_8_0, p__arg0_0_1, p___constant_11x11xf32_8_1, p__arg0_0_2, p___constant_11x11xf32_8_2, p__arg0_0_3, p___constant_11x11xf32_8_3, p__arg0_0_4, p___constant_11x11xf32_8_4, p__arg0_0_5, p___constant_11x11xf32_8_5, p__arg0_0_6, p___constant_11x11xf32_8_6, p__arg0_0_7, p___constant_11x11xf32_8_7, p__arg0_0_8, p___constant_11x11xf32_8_8, p__arg0_0_9, p___constant_11x11xf32_8_9, p__arg0_0_10, p___constant_11x11xf32_8_10) {  pe = "(0, 0, 0, 0, 8)", opr = "fmac", op_id = "17", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 start
	if (1'b1 == current_fsm_state01) begin
	    fmul_0_0_0_0_8_x <= p__arg0_0_0;
	    fmul_0_0_0_0_8_y <= p___constant_11x11xf32_8_0;
	end
	if (1'b1 == current_fsm_state03) begin
	    fadd_0_0_0_0_8_x <= p_val_cst_0_point_0000000000000000000000000;
	    fadd_0_0_0_0_8_y <= fmul_0_0_0_0_8_r;
	end

	if (1'b1 == current_fsm_state04) begin
	    fmul_0_0_0_0_8_x <= p__arg0_0_1;
	    fmul_0_0_0_0_8_y <= p___constant_11x11xf32_8_1;
	end
	if (1'b1 == current_fsm_state06) begin
	    fadd_0_0_0_0_8_x <= fadd_0_0_0_0_8_r;
	    fadd_0_0_0_0_8_y <= fmul_0_0_0_0_8_r;
	end

	if (1'b1 == current_fsm_state07) begin
	    fmul_0_0_0_0_8_x <= p__arg0_0_2;
	    fmul_0_0_0_0_8_y <= p___constant_11x11xf32_8_2;
	end
	if (1'b1 == current_fsm_state09) begin
	    fadd_0_0_0_0_8_x <= fadd_0_0_0_0_8_r;
	    fadd_0_0_0_0_8_y <= fmul_0_0_0_0_8_r;
	end

	if (1'b1 == current_fsm_state10) begin
	    fmul_0_0_0_0_8_x <= p__arg0_0_3;
	    fmul_0_0_0_0_8_y <= p___constant_11x11xf32_8_3;
	end
	if (1'b1 == current_fsm_state12) begin
	    fadd_0_0_0_0_8_x <= fadd_0_0_0_0_8_r;
	    fadd_0_0_0_0_8_y <= fmul_0_0_0_0_8_r;
	end

	if (1'b1 == current_fsm_state13) begin
	    fmul_0_0_0_0_8_x <= p__arg0_0_4;
	    fmul_0_0_0_0_8_y <= p___constant_11x11xf32_8_4;
	end
	if (1'b1 == current_fsm_state15) begin
	    fadd_0_0_0_0_8_x <= fadd_0_0_0_0_8_r;
	    fadd_0_0_0_0_8_y <= fmul_0_0_0_0_8_r;
	end

	if (1'b1 == current_fsm_state16) begin
	    fmul_0_0_0_0_8_x <= p__arg0_0_5;
	    fmul_0_0_0_0_8_y <= p___constant_11x11xf32_8_5;
	end
	if (1'b1 == current_fsm_state18) begin
	    fadd_0_0_0_0_8_x <= fadd_0_0_0_0_8_r;
	    fadd_0_0_0_0_8_y <= fmul_0_0_0_0_8_r;
	end

	if (1'b1 == current_fsm_state19) begin
	    fmul_0_0_0_0_8_x <= p__arg0_0_6;
	    fmul_0_0_0_0_8_y <= p___constant_11x11xf32_8_6;
	end
	if (1'b1 == current_fsm_state21) begin
	    fadd_0_0_0_0_8_x <= fadd_0_0_0_0_8_r;
	    fadd_0_0_0_0_8_y <= fmul_0_0_0_0_8_r;
	end

	if (1'b1 == current_fsm_state22) begin
	    fmul_0_0_0_0_8_x <= p__arg0_0_7;
	    fmul_0_0_0_0_8_y <= p___constant_11x11xf32_8_7;
	end
	if (1'b1 == current_fsm_state24) begin
	    fadd_0_0_0_0_8_x <= fadd_0_0_0_0_8_r;
	    fadd_0_0_0_0_8_y <= fmul_0_0_0_0_8_r;
	end

	if (1'b1 == current_fsm_state25) begin
	    fmul_0_0_0_0_8_x <= p__arg0_0_8;
	    fmul_0_0_0_0_8_y <= p___constant_11x11xf32_8_8;
	end
	if (1'b1 == current_fsm_state27) begin
	    fadd_0_0_0_0_8_x <= fadd_0_0_0_0_8_r;
	    fadd_0_0_0_0_8_y <= fmul_0_0_0_0_8_r;
	end

	if (1'b1 == current_fsm_state28) begin
	    fmul_0_0_0_0_8_x <= p__arg0_0_9;
	    fmul_0_0_0_0_8_y <= p___constant_11x11xf32_8_9;
	end
	if (1'b1 == current_fsm_state30) begin
	    fadd_0_0_0_0_8_x <= fadd_0_0_0_0_8_r;
	    fadd_0_0_0_0_8_y <= fmul_0_0_0_0_8_r;
	end

	if (1'b1 == current_fsm_state31) begin
	    fmul_0_0_0_0_8_x <= p__arg0_0_10;
	    fmul_0_0_0_0_8_y <= p___constant_11x11xf32_8_10;
	end
	if (1'b1 == current_fsm_state33) begin
	    fadd_0_0_0_0_8_x <= fadd_0_0_0_0_8_r;
	    fadd_0_0_0_0_8_y <= fmul_0_0_0_0_8_r;
	end

	// p_val_226 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_8_0, p__arg0_0_1, p___constant_11x11xf32_8_1, p__arg0_0_2, p___constant_11x11xf32_8_2, p__arg0_0_3, p___constant_11x11xf32_8_3, p__arg0_0_4, p___constant_11x11xf32_8_4, p__arg0_0_5, p___constant_11x11xf32_8_5, p__arg0_0_6, p___constant_11x11xf32_8_6, p__arg0_0_7, p___constant_11x11xf32_8_7, p__arg0_0_8, p___constant_11x11xf32_8_8, p__arg0_0_9, p___constant_11x11xf32_8_9, p__arg0_0_10, p___constant_11x11xf32_8_10) {  pe = "(0, 0, 0, 0, 8)", opr = "fmac", op_id = "17", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 end


	// p_val_227 = "copy" (p_val_226) {  pe = "(0, 0, 0, 0, 8)", opr = "copy", op_id = "18", start_time = "36"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state36) begin
	    p_val_227 <= fadd_0_0_0_0_8_r;
	end
	// p_val_227 = "copy" (p_val_226) {  pe = "(0, 0, 0, 0, 8)", opr = "copy", op_id = "18", start_time = "36"  } : (f32) -> f32 end


	// p_val_284 = "fadd" (p_val_227, p___constant_11xf32_8) {  pe = "(0, 0, 0, 0, 8)", opr = "fadd", op_id = "31", start_time = "37"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state37) begin
	    fadd_0_0_0_0_8_x <= p_val_227;
	    fadd_0_0_0_0_8_y <= p___constant_11xf32_8;
	end
	// p_val_284 = "fadd" (p_val_227, p___constant_11xf32_8) {  pe = "(0, 0, 0, 0, 8)", opr = "fadd", op_id = "31", start_time = "37"  } : (f32, f32) -> f32 end


	// p_val_295 = "copy" (p_val_284) {  pe = "(0, 0, 0, 0, 8)", opr = "copy", op_id = "42", start_time = "40"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state40) begin
	    p_val_295 <= fadd_0_0_0_0_8_r;
	end
	// p_val_295 = "copy" (p_val_284) {  pe = "(0, 0, 0, 0, 8)", opr = "copy", op_id = "42", start_time = "40"  } : (f32) -> f32 end


	// p_val_306 = "fadd" (p_val_295, p_val_296) {  pe = "(0, 0, 0, 0, 8)", opr = "fadd", op_id = "52", start_time = "41"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state41) begin
	    fadd_0_0_0_0_8_x <= p_val_295;
	    fadd_0_0_0_0_8_y <= p_val_296;
	end
	// p_val_306 = "fadd" (p_val_295, p_val_296) {  pe = "(0, 0, 0, 0, 8)", opr = "fadd", op_id = "52", start_time = "41"  } : (f32, f32) -> f32 end


	// p_val_307 = "copy" (p_val_297) {  pe = "(0, 0, 0, 0, 8)", opr = "copy", op_id = "53", start_time = "41"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state41) begin
	    p_val_307 <= p_val_297;
	end
	// p_val_307 = "copy" (p_val_297) {  pe = "(0, 0, 0, 0, 8)", opr = "copy", op_id = "53", start_time = "41"  } : (f32) -> f32 end


	// p_val_308 = "copy" (p_val_306) {  pe = "(0, 0, 0, 0, 8)", opr = "copy", op_id = "54", start_time = "44"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state44) begin
	    p_val_308 <= fadd_0_0_0_0_8_r;
	end
	// p_val_308 = "copy" (p_val_306) {  pe = "(0, 0, 0, 0, 8)", opr = "copy", op_id = "54", start_time = "44"  } : (f32) -> f32 end


	// p_val_309 = "fadd" (p_val_308, p_val_307) {  pe = "(0, 0, 0, 0, 8)", opr = "fadd", op_id = "55", start_time = "46"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state46) begin
	    fadd_0_0_0_0_8_x <= p_val_308;
	    fadd_0_0_0_0_8_y <= p_val_307;
	end
	// p_val_309 = "fadd" (p_val_308, p_val_307) {  pe = "(0, 0, 0, 0, 8)", opr = "fadd", op_id = "55", start_time = "46"  } : (f32, f32) -> f32 end


	// p_val_310 = "copy" (p_val_309) {  pe = "(0, 0, 0, 0, 8)", opr = "copy", op_id = "56", start_time = "49"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state49) begin
	    p_val_310 <= fadd_0_0_0_0_8_r;
	end
	// p_val_310 = "copy" (p_val_309) {  pe = "(0, 0, 0, 0, 8)", opr = "copy", op_id = "56", start_time = "49"  } : (f32) -> f32 end


	// p_val_311 = "copy" (p_val_305) {  pe = "(0, 0, 0, 0, 8)", opr = "copy", op_id = "57", start_time = "50"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state50) begin
	    p_val_311 <= fadd_0_0_0_0_0_r;
	end
	// p_val_311 = "copy" (p_val_305) {  pe = "(0, 0, 0, 0, 8)", opr = "copy", op_id = "57", start_time = "50"  } : (f32) -> f32 end


	// p_val_312 = "fadd" (p_val_311, p_val_310) {  pe = "(0, 0, 0, 0, 8)", opr = "fadd", op_id = "58", start_time = "51"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state51) begin
	    fadd_0_0_0_0_8_x <= p_val_311;
	    fadd_0_0_0_0_8_y <= p_val_310;
	end
	// p_val_312 = "fadd" (p_val_311, p_val_310) {  pe = "(0, 0, 0, 0, 8)", opr = "fadd", op_id = "58", start_time = "51"  } : (f32, f32) -> f32 end


	// p_val_313 = "copy" (p_val_312) {  pe = "(0, 0, 0, 0, 8)", opr = "copy", op_id = "59", start_time = "54"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state54) begin
	    p_val_313 <= fadd_0_0_0_0_8_r;
	end
	// p_val_313 = "copy" (p_val_312) {  pe = "(0, 0, 0, 0, 8)", opr = "copy", op_id = "59", start_time = "54"  } : (f32) -> f32 end

end

always @ (posedge clk) begin

	// p_val_250 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_9_0, p__arg0_0_1, p___constant_11x11xf32_9_1, p__arg0_0_2, p___constant_11x11xf32_9_2, p__arg0_0_3, p___constant_11x11xf32_9_3, p__arg0_0_4, p___constant_11x11xf32_9_4, p__arg0_0_5, p___constant_11x11xf32_9_5, p__arg0_0_6, p___constant_11x11xf32_9_6, p__arg0_0_7, p___constant_11x11xf32_9_7, p__arg0_0_8, p___constant_11x11xf32_9_8, p__arg0_0_9, p___constant_11x11xf32_9_9, p__arg0_0_10, p___constant_11x11xf32_9_10) {  pe = "(0, 0, 0, 0, 9)", opr = "fmac", op_id = "19", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 start
	if (1'b1 == current_fsm_state01) begin
	    fmul_0_0_0_0_9_x <= p__arg0_0_0;
	    fmul_0_0_0_0_9_y <= p___constant_11x11xf32_9_0;
	end
	if (1'b1 == current_fsm_state03) begin
	    fadd_0_0_0_0_9_x <= p_val_cst_0_point_0000000000000000000000000;
	    fadd_0_0_0_0_9_y <= fmul_0_0_0_0_9_r;
	end

	if (1'b1 == current_fsm_state04) begin
	    fmul_0_0_0_0_9_x <= p__arg0_0_1;
	    fmul_0_0_0_0_9_y <= p___constant_11x11xf32_9_1;
	end
	if (1'b1 == current_fsm_state06) begin
	    fadd_0_0_0_0_9_x <= fadd_0_0_0_0_9_r;
	    fadd_0_0_0_0_9_y <= fmul_0_0_0_0_9_r;
	end

	if (1'b1 == current_fsm_state07) begin
	    fmul_0_0_0_0_9_x <= p__arg0_0_2;
	    fmul_0_0_0_0_9_y <= p___constant_11x11xf32_9_2;
	end
	if (1'b1 == current_fsm_state09) begin
	    fadd_0_0_0_0_9_x <= fadd_0_0_0_0_9_r;
	    fadd_0_0_0_0_9_y <= fmul_0_0_0_0_9_r;
	end

	if (1'b1 == current_fsm_state10) begin
	    fmul_0_0_0_0_9_x <= p__arg0_0_3;
	    fmul_0_0_0_0_9_y <= p___constant_11x11xf32_9_3;
	end
	if (1'b1 == current_fsm_state12) begin
	    fadd_0_0_0_0_9_x <= fadd_0_0_0_0_9_r;
	    fadd_0_0_0_0_9_y <= fmul_0_0_0_0_9_r;
	end

	if (1'b1 == current_fsm_state13) begin
	    fmul_0_0_0_0_9_x <= p__arg0_0_4;
	    fmul_0_0_0_0_9_y <= p___constant_11x11xf32_9_4;
	end
	if (1'b1 == current_fsm_state15) begin
	    fadd_0_0_0_0_9_x <= fadd_0_0_0_0_9_r;
	    fadd_0_0_0_0_9_y <= fmul_0_0_0_0_9_r;
	end

	if (1'b1 == current_fsm_state16) begin
	    fmul_0_0_0_0_9_x <= p__arg0_0_5;
	    fmul_0_0_0_0_9_y <= p___constant_11x11xf32_9_5;
	end
	if (1'b1 == current_fsm_state18) begin
	    fadd_0_0_0_0_9_x <= fadd_0_0_0_0_9_r;
	    fadd_0_0_0_0_9_y <= fmul_0_0_0_0_9_r;
	end

	if (1'b1 == current_fsm_state19) begin
	    fmul_0_0_0_0_9_x <= p__arg0_0_6;
	    fmul_0_0_0_0_9_y <= p___constant_11x11xf32_9_6;
	end
	if (1'b1 == current_fsm_state21) begin
	    fadd_0_0_0_0_9_x <= fadd_0_0_0_0_9_r;
	    fadd_0_0_0_0_9_y <= fmul_0_0_0_0_9_r;
	end

	if (1'b1 == current_fsm_state22) begin
	    fmul_0_0_0_0_9_x <= p__arg0_0_7;
	    fmul_0_0_0_0_9_y <= p___constant_11x11xf32_9_7;
	end
	if (1'b1 == current_fsm_state24) begin
	    fadd_0_0_0_0_9_x <= fadd_0_0_0_0_9_r;
	    fadd_0_0_0_0_9_y <= fmul_0_0_0_0_9_r;
	end

	if (1'b1 == current_fsm_state25) begin
	    fmul_0_0_0_0_9_x <= p__arg0_0_8;
	    fmul_0_0_0_0_9_y <= p___constant_11x11xf32_9_8;
	end
	if (1'b1 == current_fsm_state27) begin
	    fadd_0_0_0_0_9_x <= fadd_0_0_0_0_9_r;
	    fadd_0_0_0_0_9_y <= fmul_0_0_0_0_9_r;
	end

	if (1'b1 == current_fsm_state28) begin
	    fmul_0_0_0_0_9_x <= p__arg0_0_9;
	    fmul_0_0_0_0_9_y <= p___constant_11x11xf32_9_9;
	end
	if (1'b1 == current_fsm_state30) begin
	    fadd_0_0_0_0_9_x <= fadd_0_0_0_0_9_r;
	    fadd_0_0_0_0_9_y <= fmul_0_0_0_0_9_r;
	end

	if (1'b1 == current_fsm_state31) begin
	    fmul_0_0_0_0_9_x <= p__arg0_0_10;
	    fmul_0_0_0_0_9_y <= p___constant_11x11xf32_9_10;
	end
	if (1'b1 == current_fsm_state33) begin
	    fadd_0_0_0_0_9_x <= fadd_0_0_0_0_9_r;
	    fadd_0_0_0_0_9_y <= fmul_0_0_0_0_9_r;
	end

	// p_val_250 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_9_0, p__arg0_0_1, p___constant_11x11xf32_9_1, p__arg0_0_2, p___constant_11x11xf32_9_2, p__arg0_0_3, p___constant_11x11xf32_9_3, p__arg0_0_4, p___constant_11x11xf32_9_4, p__arg0_0_5, p___constant_11x11xf32_9_5, p__arg0_0_6, p___constant_11x11xf32_9_6, p__arg0_0_7, p___constant_11x11xf32_9_7, p__arg0_0_8, p___constant_11x11xf32_9_8, p__arg0_0_9, p___constant_11x11xf32_9_9, p__arg0_0_10, p___constant_11x11xf32_9_10) {  pe = "(0, 0, 0, 0, 9)", opr = "fmac", op_id = "19", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 end


	// p_val_251 = "copy" (p_val_250) {  pe = "(0, 0, 0, 0, 9)", opr = "copy", op_id = "20", start_time = "36"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state36) begin
	    p_val_251 <= fadd_0_0_0_0_9_r;
	end
	// p_val_251 = "copy" (p_val_250) {  pe = "(0, 0, 0, 0, 9)", opr = "copy", op_id = "20", start_time = "36"  } : (f32) -> f32 end


	// p_val_285 = "fadd" (p_val_251, p___constant_11xf32_9) {  pe = "(0, 0, 0, 0, 9)", opr = "fadd", op_id = "32", start_time = "37"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state37) begin
	    fadd_0_0_0_0_9_x <= p_val_251;
	    fadd_0_0_0_0_9_y <= p___constant_11xf32_9;
	end
	// p_val_285 = "fadd" (p_val_251, p___constant_11xf32_9) {  pe = "(0, 0, 0, 0, 9)", opr = "fadd", op_id = "32", start_time = "37"  } : (f32, f32) -> f32 end


	// p_val_296 = "copy" (p_val_285) {  pe = "(0, 0, 0, 0, 9)", opr = "copy", op_id = "43", start_time = "40"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state40) begin
	    p_val_296 <= fadd_0_0_0_0_9_r;
	end
	// p_val_296 = "copy" (p_val_285) {  pe = "(0, 0, 0, 0, 9)", opr = "copy", op_id = "43", start_time = "40"  } : (f32) -> f32 end

end

always @ (posedge clk) begin

	// p_val_274 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_10_0, p__arg0_0_1, p___constant_11x11xf32_10_1, p__arg0_0_2, p___constant_11x11xf32_10_2, p__arg0_0_3, p___constant_11x11xf32_10_3, p__arg0_0_4, p___constant_11x11xf32_10_4, p__arg0_0_5, p___constant_11x11xf32_10_5, p__arg0_0_6, p___constant_11x11xf32_10_6, p__arg0_0_7, p___constant_11x11xf32_10_7, p__arg0_0_8, p___constant_11x11xf32_10_8, p__arg0_0_9, p___constant_11x11xf32_10_9, p__arg0_0_10, p___constant_11x11xf32_10_10) {  pe = "(0, 0, 0, 0, 10)", opr = "fmac", op_id = "21", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 start
	if (1'b1 == current_fsm_state01) begin
	    fmul_0_0_0_0_10_x <= p__arg0_0_0;
	    fmul_0_0_0_0_10_y <= p___constant_11x11xf32_10_0;
	end
	if (1'b1 == current_fsm_state03) begin
	    fadd_0_0_0_0_10_x <= p_val_cst_0_point_0000000000000000000000000;
	    fadd_0_0_0_0_10_y <= fmul_0_0_0_0_10_r;
	end

	if (1'b1 == current_fsm_state04) begin
	    fmul_0_0_0_0_10_x <= p__arg0_0_1;
	    fmul_0_0_0_0_10_y <= p___constant_11x11xf32_10_1;
	end
	if (1'b1 == current_fsm_state06) begin
	    fadd_0_0_0_0_10_x <= fadd_0_0_0_0_10_r;
	    fadd_0_0_0_0_10_y <= fmul_0_0_0_0_10_r;
	end

	if (1'b1 == current_fsm_state07) begin
	    fmul_0_0_0_0_10_x <= p__arg0_0_2;
	    fmul_0_0_0_0_10_y <= p___constant_11x11xf32_10_2;
	end
	if (1'b1 == current_fsm_state09) begin
	    fadd_0_0_0_0_10_x <= fadd_0_0_0_0_10_r;
	    fadd_0_0_0_0_10_y <= fmul_0_0_0_0_10_r;
	end

	if (1'b1 == current_fsm_state10) begin
	    fmul_0_0_0_0_10_x <= p__arg0_0_3;
	    fmul_0_0_0_0_10_y <= p___constant_11x11xf32_10_3;
	end
	if (1'b1 == current_fsm_state12) begin
	    fadd_0_0_0_0_10_x <= fadd_0_0_0_0_10_r;
	    fadd_0_0_0_0_10_y <= fmul_0_0_0_0_10_r;
	end

	if (1'b1 == current_fsm_state13) begin
	    fmul_0_0_0_0_10_x <= p__arg0_0_4;
	    fmul_0_0_0_0_10_y <= p___constant_11x11xf32_10_4;
	end
	if (1'b1 == current_fsm_state15) begin
	    fadd_0_0_0_0_10_x <= fadd_0_0_0_0_10_r;
	    fadd_0_0_0_0_10_y <= fmul_0_0_0_0_10_r;
	end

	if (1'b1 == current_fsm_state16) begin
	    fmul_0_0_0_0_10_x <= p__arg0_0_5;
	    fmul_0_0_0_0_10_y <= p___constant_11x11xf32_10_5;
	end
	if (1'b1 == current_fsm_state18) begin
	    fadd_0_0_0_0_10_x <= fadd_0_0_0_0_10_r;
	    fadd_0_0_0_0_10_y <= fmul_0_0_0_0_10_r;
	end

	if (1'b1 == current_fsm_state19) begin
	    fmul_0_0_0_0_10_x <= p__arg0_0_6;
	    fmul_0_0_0_0_10_y <= p___constant_11x11xf32_10_6;
	end
	if (1'b1 == current_fsm_state21) begin
	    fadd_0_0_0_0_10_x <= fadd_0_0_0_0_10_r;
	    fadd_0_0_0_0_10_y <= fmul_0_0_0_0_10_r;
	end

	if (1'b1 == current_fsm_state22) begin
	    fmul_0_0_0_0_10_x <= p__arg0_0_7;
	    fmul_0_0_0_0_10_y <= p___constant_11x11xf32_10_7;
	end
	if (1'b1 == current_fsm_state24) begin
	    fadd_0_0_0_0_10_x <= fadd_0_0_0_0_10_r;
	    fadd_0_0_0_0_10_y <= fmul_0_0_0_0_10_r;
	end

	if (1'b1 == current_fsm_state25) begin
	    fmul_0_0_0_0_10_x <= p__arg0_0_8;
	    fmul_0_0_0_0_10_y <= p___constant_11x11xf32_10_8;
	end
	if (1'b1 == current_fsm_state27) begin
	    fadd_0_0_0_0_10_x <= fadd_0_0_0_0_10_r;
	    fadd_0_0_0_0_10_y <= fmul_0_0_0_0_10_r;
	end

	if (1'b1 == current_fsm_state28) begin
	    fmul_0_0_0_0_10_x <= p__arg0_0_9;
	    fmul_0_0_0_0_10_y <= p___constant_11x11xf32_10_9;
	end
	if (1'b1 == current_fsm_state30) begin
	    fadd_0_0_0_0_10_x <= fadd_0_0_0_0_10_r;
	    fadd_0_0_0_0_10_y <= fmul_0_0_0_0_10_r;
	end

	if (1'b1 == current_fsm_state31) begin
	    fmul_0_0_0_0_10_x <= p__arg0_0_10;
	    fmul_0_0_0_0_10_y <= p___constant_11x11xf32_10_10;
	end
	if (1'b1 == current_fsm_state33) begin
	    fadd_0_0_0_0_10_x <= fadd_0_0_0_0_10_r;
	    fadd_0_0_0_0_10_y <= fmul_0_0_0_0_10_r;
	end

	// p_val_274 = "fmac" (p_val_cst_0_point_0000000000000000000000000, p__arg0_0_0, p___constant_11x11xf32_10_0, p__arg0_0_1, p___constant_11x11xf32_10_1, p__arg0_0_2, p___constant_11x11xf32_10_2, p__arg0_0_3, p___constant_11x11xf32_10_3, p__arg0_0_4, p___constant_11x11xf32_10_4, p__arg0_0_5, p___constant_11x11xf32_10_5, p__arg0_0_6, p___constant_11x11xf32_10_6, p__arg0_0_7, p___constant_11x11xf32_10_7, p__arg0_0_8, p___constant_11x11xf32_10_8, p__arg0_0_9, p___constant_11x11xf32_10_9, p__arg0_0_10, p___constant_11x11xf32_10_10) {  pe = "(0, 0, 0, 0, 10)", opr = "fmac", op_id = "21", start_time = "1"  } : (f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32, f32) -> f32 end


	// p_val_275 = "copy" (p_val_274) {  pe = "(0, 0, 0, 0, 10)", opr = "copy", op_id = "22", start_time = "36"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state36) begin
	    p_val_275 <= fadd_0_0_0_0_10_r;
	end
	// p_val_275 = "copy" (p_val_274) {  pe = "(0, 0, 0, 0, 10)", opr = "copy", op_id = "22", start_time = "36"  } : (f32) -> f32 end


	// p_val_286 = "fadd" (p_val_275, p___constant_11xf32_10) {  pe = "(0, 0, 0, 0, 10)", opr = "fadd", op_id = "33", start_time = "37"  } : (f32, f32) -> f32 start
	if (1'b1 == current_fsm_state37) begin
	    fadd_0_0_0_0_10_x <= p_val_275;
	    fadd_0_0_0_0_10_y <= p___constant_11xf32_10;
	end
	// p_val_286 = "fadd" (p_val_275, p___constant_11xf32_10) {  pe = "(0, 0, 0, 0, 10)", opr = "fadd", op_id = "33", start_time = "37"  } : (f32, f32) -> f32 end


	// p_val_297 = "copy" (p_val_286) {  pe = "(0, 0, 0, 0, 10)", opr = "copy", op_id = "44", start_time = "40"  } : (f32) -> f32 start
	if (1'b1 == current_fsm_state40) begin
	    p_val_297 <= fadd_0_0_0_0_10_r;
	end
	// p_val_297 = "copy" (p_val_286) {  pe = "(0, 0, 0, 0, 10)", opr = "copy", op_id = "44", start_time = "40"  } : (f32) -> f32 end

end

always @ (posedge clk) begin
    if (rst == 1'b1) begin
        current_fsm <= fsm_state01;
    end else begin
        current_fsm <= next_state_fsm;
    end
end

always @ (*) begin
    case (current_fsm)
		fsm_state01 : begin
		    next_state_fsm = fsm_state02;
		end
		fsm_state02 : begin
		    next_state_fsm = fsm_state03;
		end
		fsm_state03 : begin
		    next_state_fsm = fsm_state04;
		end
		fsm_state04 : begin
		    next_state_fsm = fsm_state05;
		end
		fsm_state05 : begin
		    next_state_fsm = fsm_state06;
		end
		fsm_state06 : begin
		    next_state_fsm = fsm_state07;
		end
		fsm_state07 : begin
		    next_state_fsm = fsm_state08;
		end
		fsm_state08 : begin
		    next_state_fsm = fsm_state09;
		end
		fsm_state09 : begin
		    next_state_fsm = fsm_state10;
		end
		fsm_state10 : begin
		    next_state_fsm = fsm_state11;
		end
		fsm_state11 : begin
		    next_state_fsm = fsm_state12;
		end
		fsm_state12 : begin
		    next_state_fsm = fsm_state13;
		end
		fsm_state13 : begin
		    next_state_fsm = fsm_state14;
		end
		fsm_state14 : begin
		    next_state_fsm = fsm_state15;
		end
		fsm_state15 : begin
		    next_state_fsm = fsm_state16;
		end
		fsm_state16 : begin
		    next_state_fsm = fsm_state17;
		end
		fsm_state17 : begin
		    next_state_fsm = fsm_state18;
		end
		fsm_state18 : begin
		    next_state_fsm = fsm_state19;
		end
		fsm_state19 : begin
		    next_state_fsm = fsm_state20;
		end
		fsm_state20 : begin
		    next_state_fsm = fsm_state21;
		end
		fsm_state21 : begin
		    next_state_fsm = fsm_state22;
		end
		fsm_state22 : begin
		    next_state_fsm = fsm_state23;
		end
		fsm_state23 : begin
		    next_state_fsm = fsm_state24;
		end
		fsm_state24 : begin
		    next_state_fsm = fsm_state25;
		end
		fsm_state25 : begin
		    next_state_fsm = fsm_state26;
		end
		fsm_state26 : begin
		    next_state_fsm = fsm_state27;
		end
		fsm_state27 : begin
		    next_state_fsm = fsm_state28;
		end
		fsm_state28 : begin
		    next_state_fsm = fsm_state29;
		end
		fsm_state29 : begin
		    next_state_fsm = fsm_state30;
		end
		fsm_state30 : begin
		    next_state_fsm = fsm_state31;
		end
		fsm_state31 : begin
		    next_state_fsm = fsm_state32;
		end
		fsm_state32 : begin
		    next_state_fsm = fsm_state33;
		end
		fsm_state33 : begin
		    next_state_fsm = fsm_state34;
		end
		fsm_state34 : begin
		    next_state_fsm = fsm_state35;
		end
		fsm_state35 : begin
		    next_state_fsm = fsm_state36;
		end
		fsm_state36 : begin
		    next_state_fsm = fsm_state37;
		end
		fsm_state37 : begin
		    next_state_fsm = fsm_state38;
		end
		fsm_state38 : begin
		    next_state_fsm = fsm_state39;
		end
		fsm_state39 : begin
		    next_state_fsm = fsm_state40;
		end
		fsm_state40 : begin
		    next_state_fsm = fsm_state41;
		end
		fsm_state41 : begin
		    next_state_fsm = fsm_state42;
		end
		fsm_state42 : begin
		    next_state_fsm = fsm_state43;
		end
		fsm_state43 : begin
		    next_state_fsm = fsm_state44;
		end
		fsm_state44 : begin
		    next_state_fsm = fsm_state45;
		end
		fsm_state45 : begin
		    next_state_fsm = fsm_state46;
		end
		fsm_state46 : begin
		    next_state_fsm = fsm_state47;
		end
		fsm_state47 : begin
		    next_state_fsm = fsm_state48;
		end
		fsm_state48 : begin
		    next_state_fsm = fsm_state49;
		end
		fsm_state49 : begin
		    next_state_fsm = fsm_state50;
		end
		fsm_state50 : begin
		    next_state_fsm = fsm_state51;
		end
		fsm_state51 : begin
		    next_state_fsm = fsm_state52;
		end
		fsm_state52 : begin
		    next_state_fsm = fsm_state53;
		end
		fsm_state53 : begin
		    next_state_fsm = fsm_state54;
		end
		fsm_state54 : begin
		    next_state_fsm = fsm_state55;
		end
		fsm_state55 : begin
		    next_state_fsm = fsm_state01;
		end
		default : begin
		    next_state_fsm = 'bx;
		end
    endcase
end
assign current_fsm_state01 = current_fsm[6'd0];
assign current_fsm_state02 = current_fsm[6'd1];
assign current_fsm_state03 = current_fsm[6'd2];
assign current_fsm_state04 = current_fsm[6'd3];
assign current_fsm_state05 = current_fsm[6'd4];
assign current_fsm_state06 = current_fsm[6'd5];
assign current_fsm_state07 = current_fsm[6'd6];
assign current_fsm_state08 = current_fsm[6'd7];
assign current_fsm_state09 = current_fsm[6'd8];
assign current_fsm_state10 = current_fsm[6'd9];
assign current_fsm_state11 = current_fsm[6'd10];
assign current_fsm_state12 = current_fsm[6'd11];
assign current_fsm_state13 = current_fsm[6'd12];
assign current_fsm_state14 = current_fsm[6'd13];
assign current_fsm_state15 = current_fsm[6'd14];
assign current_fsm_state16 = current_fsm[6'd15];
assign current_fsm_state17 = current_fsm[6'd16];
assign current_fsm_state18 = current_fsm[6'd17];
assign current_fsm_state19 = current_fsm[6'd18];
assign current_fsm_state20 = current_fsm[6'd19];
assign current_fsm_state21 = current_fsm[6'd20];
assign current_fsm_state22 = current_fsm[6'd21];
assign current_fsm_state23 = current_fsm[6'd22];
assign current_fsm_state24 = current_fsm[6'd23];
assign current_fsm_state25 = current_fsm[6'd24];
assign current_fsm_state26 = current_fsm[6'd25];
assign current_fsm_state27 = current_fsm[6'd26];
assign current_fsm_state28 = current_fsm[6'd27];
assign current_fsm_state29 = current_fsm[6'd28];
assign current_fsm_state30 = current_fsm[6'd29];
assign current_fsm_state31 = current_fsm[6'd30];
assign current_fsm_state32 = current_fsm[6'd31];
assign current_fsm_state33 = current_fsm[6'd32];
assign current_fsm_state34 = current_fsm[6'd33];
assign current_fsm_state35 = current_fsm[6'd34];
assign current_fsm_state36 = current_fsm[6'd35];
assign current_fsm_state37 = current_fsm[6'd36];
assign current_fsm_state38 = current_fsm[6'd37];
assign current_fsm_state39 = current_fsm[6'd38];
assign current_fsm_state40 = current_fsm[6'd39];
assign current_fsm_state41 = current_fsm[6'd40];
assign current_fsm_state42 = current_fsm[6'd41];
assign current_fsm_state43 = current_fsm[6'd42];
assign current_fsm_state44 = current_fsm[6'd43];
assign current_fsm_state45 = current_fsm[6'd44];
assign current_fsm_state46 = current_fsm[6'd45];
assign current_fsm_state47 = current_fsm[6'd46];
assign current_fsm_state48 = current_fsm[6'd47];
assign current_fsm_state49 = current_fsm[6'd48];
assign current_fsm_state50 = current_fsm[6'd49];
assign current_fsm_state51 = current_fsm[6'd50];
assign current_fsm_state52 = current_fsm[6'd51];
assign current_fsm_state53 = current_fsm[6'd52];
assign current_fsm_state54 = current_fsm[6'd53];
assign current_fsm_state55 = current_fsm[6'd54];


assign output_p_val_313 = p_val_313;

`ifdef COCOTB_SIM
initial begin
  $dumpfile ("linear.vcd");
  $dumpvars (0, linear);
  #1;
end
`endif


endmodule

